
entity TEST_REMOTE_DIMMER is
end entity;


