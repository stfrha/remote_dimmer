-- Xilinx Vhdl produced by program ngd2vhdl C.22
-- Command: -w REMOTE_DIMMER.nga time_sim.vhd 
-- Options: -w -ti UUT 
-- Date: Thu Apr 12 13:53:17 2001 
-- Input file: REMOTE_DIMMER.nga
-- Output file: time_sim.vhd
-- Tmp file: D:/TEMP/xil_13
-- Design name: REMOTE_DIMMER
-- Xilinx: W:/Xilinx
-- # of Entities: 1
-- Device: XC95108-7-PC84

-- The output of ngd2vhdl is a simulation model. This file cannot be synthesized,
-- or used in any other manner other than simulation. This netlist uses simulation
-- primitives which may not represent the true implementation of the device, however
-- the netlist is functionally correct. Do not modify this file.

-- Model for  ROC (Reset-On-Configuration) Cell
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.VITAL_Timing.all;
entity ROC is
  generic (InstancePath: STRING := "*";
           WIDTH : Time := 100 ns);
  port(O : out std_ulogic := '1') ;
  attribute VITAL_LEVEL0 of ROC : entity is TRUE;
end ROC;

architecture ROC_V of ROC is
attribute VITAL_LEVEL0 of ROC_V : architecture is TRUE;
begin
  ONE_SHOT : process
  begin
    if (WIDTH <= 0 ns) then
       assert FALSE report
       "*** Error: a positive value of WIDTH must be specified ***"
       severity failure;
    else
       wait for WIDTH;
       O <= '0';
    end if;
    wait;
  end process ONE_SHOT;
end ROC_V;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library SIMPRIM;
use SIMPRIM.VCOMPONENTS.ALL;
use SIMPRIM.VPACKAGE.ALL;
entity REMOTE_DIMMER is 
  port (
    CLK : in STD_LOGIC := 'X'; 
    RESET : in STD_LOGIC := 'X'; 
    IR_DETECT : in STD_LOGIC := 'X'; 
    ZERO_DETECT : in STD_LOGIC := 'X'; 
    TRIAC_PULSE : out STD_LOGIC; 
    RC_ADDRESS : in STD_LOGIC_VECTOR ( 3 downto 0 ) 
  );
end REMOTE_DIMMER;

architecture STRUCTURE of REMOTE_DIMMER is
  component ROC
    generic (InstancePath: STRING := "*";
             WIDTH : Time := 100 ns);
    port (O : out STD_ULOGIC := '1');
  end component;
  signal TD1_TRIAC_TRIG_I : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_Q : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D1 : STD_LOGIC; 
  signal EXP1_EXP : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D2_PT_0 : STD_LOGIC; 
  signal TD1_CNT_5_Q_0 : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D2_PT_1 : STD_LOGIC; 
  signal LIGHT_VALUE_4_FBK : STD_LOGIC; 
  signal TD1_CNT_4_Q_1 : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D2_PT_2 : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D2_PT_3 : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_UIM : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D2_PT_4 : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D2_PT_5 : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D2 : STD_LOGIC; 
  signal EXP1_EXP_PT_0 : STD_LOGIC; 
  signal EXP1_EXP_PT_1 : STD_LOGIC; 
  signal LIGHT_VALUE_4_Q : STD_LOGIC; 
  signal LIGHT_VALUE_4_RSTF : STD_LOGIC; 
  signal LIGHT_VALUE_4_R_OR_PRLD : STD_LOGIC; 
  signal LIGHT_VALUE_4_D : STD_LOGIC; 
  signal CLK_C_FCLK : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK : STD_LOGIC; 
  signal LIGHT_VALUE_4_RSTF_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_4_D1 : STD_LOGIC; 
  signal EXP0_EXP : STD_LOGIC; 
  signal LIGHT_VALUE_4_D2_PT_0 : STD_LOGIC; 
  signal FC1_CNT_3_FBK : STD_LOGIC; 
  signal FC1_CNT_4_FBK : STD_LOGIC; 
  signal FC1_CNT_5_FBK : STD_LOGIC; 
  signal FC1_CNT_6_FBK : STD_LOGIC; 
  signal FC1_CNT_7_FBK : STD_LOGIC; 
  signal LIGHT_VALUE_4_D2_PT_1 : STD_LOGIC; 
  signal LIGHT_VALUE_4_D2 : STD_LOGIC; 
  signal LIGHT_VALUE_4_D_TFF : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_1 : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_2 : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP : STD_LOGIC; 
  signal EXP0_EXP_PT_0 : STD_LOGIC; 
  signal EXP0_EXP_PT_1 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_Q : STD_LOGIC; 
  signal FSRIO_0 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_R_OR_PRLD : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D1 : STD_LOGIC; 
  signal EXP2_EXP : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D2_PT_0 : STD_LOGIC; 
  signal CM_PANIC_ON : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D2_PT_1 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D2 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D_TFF : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_0 : STD_LOGIC; 
  signal CM_FADE_UP : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_1 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP : STD_LOGIC; 
  signal CM_FADE_DOWN : STD_LOGIC; 
  signal EXP2_EXP_PT_0 : STD_LOGIC; 
  signal EXP2_EXP_PT_1 : STD_LOGIC; 
  signal EXP2_EXP_PT_2 : STD_LOGIC; 
  signal EXP2_EXP_PT_3 : STD_LOGIC; 
  signal CM_FADE_DOWN_Q : STD_LOGIC; 
  signal CM_FADE_DOWN_R_OR_PRLD : STD_LOGIC; 
  signal CM_FADE_DOWN_D : STD_LOGIC; 
  signal CM_FADE_DOWN_D1 : STD_LOGIC; 
  signal RXD_ACK : STD_LOGIC; 
  signal CM_FADE_DOWN_D2_PT_0 : STD_LOGIC; 
  signal RXD_2_FBK : STD_LOGIC; 
  signal CM_FADE_DOWN_D2_PT_1 : STD_LOGIC; 
  signal RXD_READY_FBK : STD_LOGIC; 
  signal CM_FADE_DOWN_D2_PT_2 : STD_LOGIC; 
  signal EXP19_EXP : STD_LOGIC; 
  signal CM_FADE_DOWN_D2_PT_3 : STD_LOGIC; 
  signal EXP20_EXP : STD_LOGIC; 
  signal CM_FADE_DOWN_D2_PT_4 : STD_LOGIC; 
  signal RXD_4_FBK : STD_LOGIC; 
  signal CM_FADE_DOWN_D2_PT_5 : STD_LOGIC; 
  signal CM_FADE_DOWN_D2_PT_6 : STD_LOGIC; 
  signal CM_FADE_DOWN_D2 : STD_LOGIC; 
  signal CM_FADE_DOWN_D_TFF : STD_LOGIC; 
  signal CM_FADE_DOWN_FBK : STD_LOGIC; 
  signal RXD_ACK_Q : STD_LOGIC; 
  signal RXD_ACK_R_OR_PRLD : STD_LOGIC; 
  signal RXD_ACK_D : STD_LOGIC; 
  signal RXD_ACK_D1 : STD_LOGIC; 
  signal RXD_READY : STD_LOGIC; 
  signal RXD_ACK_D2_PT_0 : STD_LOGIC; 
  signal RXD_ACK_D2 : STD_LOGIC; 
  signal RXD_READY_Q : STD_LOGIC; 
  signal RXD_READY_R_OR_PRLD : STD_LOGIC; 
  signal RXD_READY_D : STD_LOGIC; 
  signal RXD_READY_D1 : STD_LOGIC; 
  signal RXD_7_EXP : STD_LOGIC; 
  signal RXD_READY_D2_PT_0 : STD_LOGIC; 
  signal RXD_READY_D2 : STD_LOGIC; 
  signal RXD_5_FBK : STD_LOGIC; 
  signal RXD_READY_EXP_PT_0 : STD_LOGIC; 
  signal RXD_READY_EXP_PT_1 : STD_LOGIC; 
  signal RXD_6_FBK : STD_LOGIC; 
  signal RXD_READY_EXP_PT_2 : STD_LOGIC; 
  signal RXD_READY_EXP_PT_3 : STD_LOGIC; 
  signal RXD_7_FBK : STD_LOGIC; 
  signal RXD_READY_EXP_PT_4 : STD_LOGIC; 
  signal RXD_READY_EXP : STD_LOGIC; 
  signal UAR1_BYTE_AVAIL : STD_LOGIC; 
  signal RXD_7_EXP_PT_0 : STD_LOGIC; 
  signal RXD_7_EXP_PT_1 : STD_LOGIC; 
  signal RXD_7_Q : STD_LOGIC; 
  signal RXD_7_R_OR_PRLD : STD_LOGIC; 
  signal RXD_7_D : STD_LOGIC; 
  signal RXD_7_D1 : STD_LOGIC; 
  signal RXD_7_D2_PT_0 : STD_LOGIC; 
  signal RXD_7_D2_PT_1 : STD_LOGIC; 
  signal RXD_7_D2 : STD_LOGIC; 
  signal RXD_7_D_TFF : STD_LOGIC; 
  signal UAR1_BYTE_AVAIL_Q : STD_LOGIC; 
  signal UAR1_BYTE_AVAIL_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BYTE_AVAIL_D : STD_LOGIC; 
  signal UAR1_BYTE_AVAIL_D1 : STD_LOGIC; 
  signal UAR1_BIT_DONE_FBK : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_Q_4 : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_0_FBK : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_1_FBK : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_2_FBK : STD_LOGIC; 
  signal UAR1_BYTE_AVAIL_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BYTE_AVAIL_D2 : STD_LOGIC; 
  signal UAR1_BYTE_AVAIL_FBK : STD_LOGIC; 
  signal UAR1_BIT_DONE_Q : STD_LOGIC; 
  signal UAR1_BIT_DONE : STD_LOGIC; 
  signal UAR1_BIT_DONE_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BIT_DONE_D : STD_LOGIC; 
  signal UAR1_BIT_DONE_D1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_Q_5 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_1_FBK : STD_LOGIC; 
  signal UAR1_BIT_DONE_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BIT_DONE_D2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_Q : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D1 : STD_LOGIC; 
  signal EXP9_EXP : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_0 : STD_LOGIC; 
  signal EXP10_EXP : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_FBK : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_10_Q_6 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_FBK : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_FBK : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_3 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_FBK : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_4 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_FBK : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_5 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_FBK : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_6 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2 : STD_LOGIC; 
  signal UAR1_DATA_IN : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_FBK : STD_LOGIC; 
  signal EXP9_EXP_PT_0 : STD_LOGIC; 
  signal EXP9_EXP_PT_1 : STD_LOGIC; 
  signal EXP9_EXP_PT_2 : STD_LOGIC; 
  signal EXP9_EXP_PT_3 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_FBK : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_FBK : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_9_FBK : STD_LOGIC; 
  signal EXP9_EXP_PT_4 : STD_LOGIC; 
  signal UAR1_DATA_IN_Q : STD_LOGIC; 
  signal UAR1_DATA_IN_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_DATA_IN_D : STD_LOGIC; 
  signal UAR1_DATA_IN_D1 : STD_LOGIC; 
  signal IR_DETECT_C : STD_LOGIC; 
  signal UAR1_DATA_IN_D2_PT_0 : STD_LOGIC; 
  signal UAR1_DATA_IN_D2 : STD_LOGIC; 
  signal UAR1_DATA_IN_FBK : STD_LOGIC; 
  signal RESET_C : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_0_Q : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_0_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_0_D : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_0_D1 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_3_FBK : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_0_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_0_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_0_D2 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_3_Q : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_3_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_3_D : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_3_D1 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_3_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_FBK : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_3_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_3_D2 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_Q : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D1 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_2_FBK : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_1_Q : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_1_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_1_D : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_1_D1 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_1_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_1_D2 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_2_Q : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_2_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_2_D : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_2_D1 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_2_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_2_D2 : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_1_Q : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_1_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_1_D : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_1_D1 : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_1_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_1_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_1_D2 : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_2_Q : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_2_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_2_D : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_2_D1 : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_2_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_2_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_2_D2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_Q : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_D : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_D1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_D2_PT_2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_D2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_Q : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_Q_7 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_D : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_D1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_D2_PT_2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_D2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_Q : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_Q_8 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_D : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_D1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_D2_PT_2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_D2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_Q : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_D : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_D1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_D2_PT_2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_D2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_Q : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_D : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_D1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_D2_PT_2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_D2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_Q : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_D : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_D1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_D2_PT_2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_D2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_Q : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_D : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_D1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_D2_PT_2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_D2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_Q : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_D : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_D1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_D2_PT_2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_D2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_9_Q : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_9_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_9_D : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_9_D1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_9_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_9_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_9_D2 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_10_Q : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_10_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_10_D : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_10_D1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_10_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_10_FBK : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_10_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_10_D2 : STD_LOGIC; 
  signal EXP10_EXP_PT_0 : STD_LOGIC; 
  signal EXP10_EXP_PT_1 : STD_LOGIC; 
  signal EXP10_EXP_PT_2 : STD_LOGIC; 
  signal EXP10_EXP_PT_3 : STD_LOGIC; 
  signal EXP10_EXP_PT_4 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_7_Q : STD_LOGIC; 
  signal UAR1_BYTE_OUT_7_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BYTE_OUT_7_D : STD_LOGIC; 
  signal UAR1_BYTE_OUT_7_D1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_7_FBK : STD_LOGIC; 
  signal UAR1_BYTE_OUT_7_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_7_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_7_D2 : STD_LOGIC; 
  signal RXD_5_Q : STD_LOGIC; 
  signal RXD_5_R_OR_PRLD : STD_LOGIC; 
  signal RXD_5_D : STD_LOGIC; 
  signal RXD_5_D1 : STD_LOGIC; 
  signal RXD_5_D2_PT_0 : STD_LOGIC; 
  signal RXD_5_D2_PT_1 : STD_LOGIC; 
  signal RXD_5_D2 : STD_LOGIC; 
  signal RXD_5_D_TFF : STD_LOGIC; 
  signal UAR1_BYTE_OUT_5_Q : STD_LOGIC; 
  signal UAR1_BYTE_OUT_5_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BYTE_OUT_5_D : STD_LOGIC; 
  signal UAR1_BYTE_OUT_5_D1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_5_FBK : STD_LOGIC; 
  signal UAR1_BYTE_OUT_5_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_5_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_5_D2 : STD_LOGIC; 
  signal RXD_6_Q : STD_LOGIC; 
  signal RXD_6_R_OR_PRLD : STD_LOGIC; 
  signal RXD_6_D : STD_LOGIC; 
  signal RXD_6_D1 : STD_LOGIC; 
  signal RXD_6_D2_PT_0 : STD_LOGIC; 
  signal RXD_6_D2_PT_1 : STD_LOGIC; 
  signal RXD_6_D2 : STD_LOGIC; 
  signal RXD_6_D_TFF : STD_LOGIC; 
  signal UAR1_BYTE_OUT_6_Q : STD_LOGIC; 
  signal UAR1_BYTE_OUT_6_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BYTE_OUT_6_D : STD_LOGIC; 
  signal UAR1_BYTE_OUT_6_D1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_6_FBK : STD_LOGIC; 
  signal UAR1_BYTE_OUT_6_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_6_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_6_D2 : STD_LOGIC; 
  signal RXD_2_Q : STD_LOGIC; 
  signal RXD_2_R_OR_PRLD : STD_LOGIC; 
  signal RXD_2_D : STD_LOGIC; 
  signal RXD_2_D1 : STD_LOGIC; 
  signal RXD_2_D2_PT_0 : STD_LOGIC; 
  signal RXD_2_D2_PT_1 : STD_LOGIC; 
  signal RXD_2_D2 : STD_LOGIC; 
  signal RXD_2_D_TFF : STD_LOGIC; 
  signal UAR1_BYTE_OUT_2_Q : STD_LOGIC; 
  signal UAR1_BYTE_OUT_2_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BYTE_OUT_2_D : STD_LOGIC; 
  signal UAR1_BYTE_OUT_2_D1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_2_FBK : STD_LOGIC; 
  signal UAR1_BYTE_OUT_2_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_2_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_2_D2 : STD_LOGIC; 
  signal EXP19_EXP_PT_0 : STD_LOGIC; 
  signal EXP19_EXP_PT_1 : STD_LOGIC; 
  signal EXP19_EXP_PT_2 : STD_LOGIC; 
  signal EXP19_EXP_PT_3 : STD_LOGIC; 
  signal EXP19_EXP_PT_4 : STD_LOGIC; 
  signal RXD_1_EXP : STD_LOGIC; 
  signal EXP20_EXP_PT_0 : STD_LOGIC; 
  signal RXD_3_FBK : STD_LOGIC; 
  signal EXP20_EXP_PT_1 : STD_LOGIC; 
  signal RXD_0_FBK : STD_LOGIC; 
  signal EXP20_EXP_PT_2 : STD_LOGIC; 
  signal RXD_1_FBK : STD_LOGIC; 
  signal EXP20_EXP_PT_3 : STD_LOGIC; 
  signal EXP20_EXP_PT_4 : STD_LOGIC; 
  signal EXP20_EXP_PT_5 : STD_LOGIC; 
  signal RXD_1_EXP_PT_0 : STD_LOGIC; 
  signal RXD_1_EXP_PT_1 : STD_LOGIC; 
  signal RXD_1_Q : STD_LOGIC; 
  signal RXD_1_R_OR_PRLD : STD_LOGIC; 
  signal RXD_1_D : STD_LOGIC; 
  signal RXD_1_D1 : STD_LOGIC; 
  signal RXD_1_D2_PT_0 : STD_LOGIC; 
  signal RXD_1_D2_PT_1 : STD_LOGIC; 
  signal RXD_1_D2 : STD_LOGIC; 
  signal RXD_1_D_TFF : STD_LOGIC; 
  signal UAR1_BYTE_OUT_1_Q : STD_LOGIC; 
  signal UAR1_BYTE_OUT_1_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BYTE_OUT_1_D : STD_LOGIC; 
  signal UAR1_BYTE_OUT_1_D1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_1_FBK : STD_LOGIC; 
  signal UAR1_BYTE_OUT_1_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_1_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_1_D2 : STD_LOGIC; 
  signal RXD_3_Q : STD_LOGIC; 
  signal RXD_3_R_OR_PRLD : STD_LOGIC; 
  signal RXD_3_D : STD_LOGIC; 
  signal RXD_3_D1 : STD_LOGIC; 
  signal RXD_3_D2_PT_0 : STD_LOGIC; 
  signal RXD_3_D2_PT_1 : STD_LOGIC; 
  signal RXD_3_D2 : STD_LOGIC; 
  signal RXD_3_D_TFF : STD_LOGIC; 
  signal UAR1_BYTE_OUT_3_Q : STD_LOGIC; 
  signal UAR1_BYTE_OUT_3_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BYTE_OUT_3_D : STD_LOGIC; 
  signal UAR1_BYTE_OUT_3_D1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_3_FBK : STD_LOGIC; 
  signal UAR1_BYTE_OUT_3_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_3_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_3_D2 : STD_LOGIC; 
  signal RXD_0_EXP_PT_0 : STD_LOGIC; 
  signal CM_PANIC_ON_FBK : STD_LOGIC; 
  signal RXD_0_EXP_PT_1 : STD_LOGIC; 
  signal RXD_0_EXP : STD_LOGIC; 
  signal RXD_0_Q : STD_LOGIC; 
  signal RXD_0_R_OR_PRLD : STD_LOGIC; 
  signal RXD_0_D : STD_LOGIC; 
  signal RXD_0_D1 : STD_LOGIC; 
  signal RXD_0_D2_PT_0 : STD_LOGIC; 
  signal RXD_0_D2_PT_1 : STD_LOGIC; 
  signal RXD_0_D2 : STD_LOGIC; 
  signal RXD_0_D_TFF : STD_LOGIC; 
  signal UAR1_BYTE_OUT_0_Q : STD_LOGIC; 
  signal UAR1_BYTE_OUT_0_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BYTE_OUT_0_D : STD_LOGIC; 
  signal UAR1_BYTE_OUT_0_D1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_0_FBK : STD_LOGIC; 
  signal UAR1_BYTE_OUT_0_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_0_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_0_D2 : STD_LOGIC; 
  signal CM_PANIC_ON_Q : STD_LOGIC; 
  signal CM_PANIC_ON_R_OR_PRLD : STD_LOGIC; 
  signal CM_PANIC_ON_D : STD_LOGIC; 
  signal CM_PANIC_ON_D1 : STD_LOGIC; 
  signal CM_PANIC_ON_D2_PT_0 : STD_LOGIC; 
  signal CM_PANIC_ON_D2_PT_1 : STD_LOGIC; 
  signal EXP17_EXP : STD_LOGIC; 
  signal CM_PANIC_ON_D2_PT_2 : STD_LOGIC; 
  signal EXP18_EXP : STD_LOGIC; 
  signal CM_PANIC_ON_D2_PT_3 : STD_LOGIC; 
  signal CM_PANIC_ON_D2_PT_4 : STD_LOGIC; 
  signal CM_PANIC_ON_D2_PT_5 : STD_LOGIC; 
  signal CM_PANIC_ON_D2_PT_6 : STD_LOGIC; 
  signal CM_PANIC_ON_D2 : STD_LOGIC; 
  signal CM_PANIC_ON_D_TFF : STD_LOGIC; 
  signal EXP17_EXP_PT_0 : STD_LOGIC; 
  signal EXP17_EXP_PT_1 : STD_LOGIC; 
  signal EXP17_EXP_PT_2 : STD_LOGIC; 
  signal EXP17_EXP_PT_3 : STD_LOGIC; 
  signal EXP17_EXP_PT_4 : STD_LOGIC; 
  signal EXP18_EXP_PT_0 : STD_LOGIC; 
  signal EXP18_EXP_PT_1 : STD_LOGIC; 
  signal EXP18_EXP_PT_2 : STD_LOGIC; 
  signal EXP18_EXP_PT_3 : STD_LOGIC; 
  signal EXP18_EXP_PT_4 : STD_LOGIC; 
  signal EXP18_EXP_PT_5 : STD_LOGIC; 
  signal RXD_4_Q : STD_LOGIC; 
  signal RXD_4_R_OR_PRLD : STD_LOGIC; 
  signal RXD_4_D : STD_LOGIC; 
  signal RXD_4_D1 : STD_LOGIC; 
  signal RXD_4_D2_PT_0 : STD_LOGIC; 
  signal RXD_4_D2_PT_1 : STD_LOGIC; 
  signal RXD_4_D2 : STD_LOGIC; 
  signal RXD_4_D_TFF : STD_LOGIC; 
  signal UAR1_BYTE_OUT_4_Q : STD_LOGIC; 
  signal UAR1_BYTE_OUT_4_R_OR_PRLD : STD_LOGIC; 
  signal UAR1_BYTE_OUT_4_D : STD_LOGIC; 
  signal UAR1_BYTE_OUT_4_D1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_4_FBK : STD_LOGIC; 
  signal UAR1_BYTE_OUT_4_D2_PT_0 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_4_D2_PT_1 : STD_LOGIC; 
  signal UAR1_BYTE_OUT_4_D2 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_Q : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_R_OR_PRLD : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D1 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_0 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_1 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D_TFF : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3 : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP : STD_LOGIC; 
  signal FC1_CNT_3_Q : STD_LOGIC; 
  signal FC1_CNT_3_RSTF : STD_LOGIC; 
  signal FC1_CNT_3_R_OR_PRLD : STD_LOGIC; 
  signal FC1_CNT_3_D : STD_LOGIC; 
  signal FC1_CNT_3_RSTF_PT_0 : STD_LOGIC; 
  signal FC1_CNT_3_D1 : STD_LOGIC; 
  signal EXP4_EXP : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_0 : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_1 : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2 : STD_LOGIC; 
  signal FC1_CNT_3_D2 : STD_LOGIC; 
  signal FC1_CNT_3_D_TFF : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_0 : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_1 : STD_LOGIC; 
  signal FC1_CNT_3_EXP : STD_LOGIC; 
  signal FC1_CNT_7_EXP : STD_LOGIC; 
  signal EXP4_EXP_PT_0 : STD_LOGIC; 
  signal EXP4_EXP_PT_1 : STD_LOGIC; 
  signal EXP4_EXP_PT_2 : STD_LOGIC; 
  signal EXP4_EXP_PT_3 : STD_LOGIC; 
  signal EXP4_EXP_PT_4 : STD_LOGIC; 
  signal EXP4_EXP_PT_5 : STD_LOGIC; 
  signal FC1_CNT_7_Q : STD_LOGIC; 
  signal FC1_CNT_7_RSTF : STD_LOGIC; 
  signal FC1_CNT_7_R_OR_PRLD : STD_LOGIC; 
  signal FC1_CNT_7_D : STD_LOGIC; 
  signal FC1_CNT_7_RSTF_PT_0 : STD_LOGIC; 
  signal FC1_CNT_7_D1 : STD_LOGIC; 
  signal EXP3_EXP : STD_LOGIC; 
  signal FC1_CNT_7_D2_PT_0 : STD_LOGIC; 
  signal FC1_CNT_7_D2_PT_1 : STD_LOGIC; 
  signal FC1_CNT_7_D2 : STD_LOGIC; 
  signal FC1_CNT_7_D_TFF : STD_LOGIC; 
  signal FC1_CNT_7_EXP_PT_0 : STD_LOGIC; 
  signal FC1_CNT_7_EXP_PT_1 : STD_LOGIC; 
  signal FC1_CNT_7_EXP_PT_2 : STD_LOGIC; 
  signal EXP3_EXP_PT_0 : STD_LOGIC; 
  signal EXP3_EXP_PT_1 : STD_LOGIC; 
  signal EXP3_EXP_PT_2 : STD_LOGIC; 
  signal EXP3_EXP_PT_3 : STD_LOGIC; 
  signal EXP3_EXP_PT_4 : STD_LOGIC; 
  signal EXP3_EXP_PT_5 : STD_LOGIC; 
  signal FC1_CNT_1_Q : STD_LOGIC; 
  signal FC1_CNT_1_RSTF : STD_LOGIC; 
  signal FC1_CNT_1_R_OR_PRLD : STD_LOGIC; 
  signal FC1_CNT_1_D : STD_LOGIC; 
  signal FC1_CNT_1_RSTF_PT_0 : STD_LOGIC; 
  signal FC1_CNT_1_D1 : STD_LOGIC; 
  signal FC1_CNT_0_EXP : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_5_FBK : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_1 : STD_LOGIC; 
  signal LIGHT_VALUE_1_FBK : STD_LOGIC; 
  signal LIGHT_VALUE_3_FBK : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_2 : STD_LOGIC; 
  signal LIGHT_VALUE_2_FBK : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_3 : STD_LOGIC; 
  signal FC1_CNT_1_FBK : STD_LOGIC; 
  signal FC1_CNT_2_FBK : STD_LOGIC; 
  signal LIGHT_VALUE_0_FBK : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4 : STD_LOGIC; 
  signal FC1_CNT_1_D2 : STD_LOGIC; 
  signal FC1_CNT_1_D_TFF : STD_LOGIC; 
  signal FC1_CNT_0_Q : STD_LOGIC; 
  signal FC1_CNT_0_RSTF : STD_LOGIC; 
  signal FC1_CNT_0_R_OR_PRLD : STD_LOGIC; 
  signal FC1_CNT_0_D : STD_LOGIC; 
  signal FC1_CNT_0_RSTF_PT_0 : STD_LOGIC; 
  signal FC1_CNT_0_D1 : STD_LOGIC; 
  signal EXP12_EXP : STD_LOGIC; 
  signal FC1_CNT_0_D2_PT_0 : STD_LOGIC; 
  signal FC1_CNT_0_D2_PT_1 : STD_LOGIC; 
  signal FC1_CNT_0_D2 : STD_LOGIC; 
  signal FC1_CNT_0_D_TFF : STD_LOGIC; 
  signal FC1_CNT_0_EXP_PT_0 : STD_LOGIC; 
  signal FC1_CNT_0_FBK : STD_LOGIC; 
  signal FC1_CNT_0_EXP_PT_1 : STD_LOGIC; 
  signal FC1_CNT_0_EXP_PT_2 : STD_LOGIC; 
  signal EXP12_EXP_PT_0 : STD_LOGIC; 
  signal EXP12_EXP_PT_1 : STD_LOGIC; 
  signal EXP12_EXP_PT_2 : STD_LOGIC; 
  signal EXP12_EXP_PT_3 : STD_LOGIC; 
  signal EXP12_EXP_PT_4 : STD_LOGIC; 
  signal LIGHT_VALUE_5_Q : STD_LOGIC; 
  signal LIGHT_VALUE_5_D : STD_LOGIC; 
  signal LIGHT_VALUE_5_SETF : STD_LOGIC; 
  signal LIGHT_VALUE_5_SETF_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_5_D1 : STD_LOGIC; 
  signal TD1_CNT_0_EXP : STD_LOGIC; 
  signal LIGHT_VALUE_5_D2_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_5_D2_PT_1 : STD_LOGIC; 
  signal LIGHT_VALUE_5_D2 : STD_LOGIC; 
  signal LIGHT_VALUE_5_D_TFF : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1 : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_2 : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP : STD_LOGIC; 
  signal TD1_CNT_0_Q : STD_LOGIC; 
  signal TD1_CNT_0_Q_2 : STD_LOGIC; 
  signal TD1_CNT_0_RSTF : STD_LOGIC; 
  signal TD1_CNT_0_R_OR_PRLD : STD_LOGIC; 
  signal TD1_CNT_0_D : STD_LOGIC; 
  signal TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM : STD_LOGIC; 
  signal TD1_CNT_0_RSTF_PT_0 : STD_LOGIC; 
  signal TD1_CNT_0_D1 : STD_LOGIC; 
  signal TD1_CNT_0_FBK : STD_LOGIC; 
  signal TD1_CNT_0_D2_PT_0 : STD_LOGIC; 
  signal TD1_CNT_0_D2 : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0 : STD_LOGIC; 
  signal TD1_CNT_5_TD1_CNT_5_SETF_INT_Q : STD_LOGIC; 
  signal TD1_CNT_5_TD1_CNT_5_SETF_INT_D : STD_LOGIC; 
  signal TD1_CNT_5_TD1_CNT_5_SETF_INT_D1 : STD_LOGIC; 
  signal ZERO_DETECT_C : STD_LOGIC; 
  signal TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0 : STD_LOGIC; 
  signal TD1_CNT_5_TD1_CNT_5_SETF_INT_D2 : STD_LOGIC; 
  signal TD1_CNT_5_TD1_CNT_5_SETF_INT_FBK : STD_LOGIC; 
  signal FC1_CNT_2_Q : STD_LOGIC; 
  signal FC1_CNT_2_RSTF : STD_LOGIC; 
  signal FC1_CNT_2_R_OR_PRLD : STD_LOGIC; 
  signal FC1_CNT_2_D : STD_LOGIC; 
  signal FC1_CNT_2_RSTF_PT_0 : STD_LOGIC; 
  signal FC1_CNT_2_D1 : STD_LOGIC; 
  signal EXP14_EXP : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_0 : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_1 : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2 : STD_LOGIC; 
  signal FC1_CNT_2_D2 : STD_LOGIC; 
  signal FC1_CNT_2_D_TFF : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_0 : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_1 : STD_LOGIC; 
  signal FC1_CNT_2_EXP : STD_LOGIC; 
  signal LIGHT_VALUE_1_EXP : STD_LOGIC; 
  signal EXP14_EXP_PT_0 : STD_LOGIC; 
  signal EXP14_EXP_PT_1 : STD_LOGIC; 
  signal EXP14_EXP_PT_2 : STD_LOGIC; 
  signal EXP14_EXP_PT_3 : STD_LOGIC; 
  signal EXP14_EXP_PT_4 : STD_LOGIC; 
  signal EXP14_EXP_PT_5 : STD_LOGIC; 
  signal LIGHT_VALUE_1_Q : STD_LOGIC; 
  signal LIGHT_VALUE_1_D : STD_LOGIC; 
  signal LIGHT_VALUE_1_SETF : STD_LOGIC; 
  signal LIGHT_VALUE_1_SETF_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_1_D1 : STD_LOGIC; 
  signal EXP13_EXP : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_1 : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_2 : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_3 : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2 : STD_LOGIC; 
  signal LIGHT_VALUE_1_D_TFF : STD_LOGIC; 
  signal LIGHT_VALUE_1_EXP_PT_0 : STD_LOGIC; 
  signal EXP13_EXP_PT_0 : STD_LOGIC; 
  signal EXP13_EXP_PT_1 : STD_LOGIC; 
  signal EXP13_EXP_PT_2 : STD_LOGIC; 
  signal EXP13_EXP_PT_3 : STD_LOGIC; 
  signal EXP13_EXP_PT_4 : STD_LOGIC; 
  signal FC1_CNT_4_Q : STD_LOGIC; 
  signal FC1_CNT_4_RSTF : STD_LOGIC; 
  signal FC1_CNT_4_R_OR_PRLD : STD_LOGIC; 
  signal FC1_CNT_4_D : STD_LOGIC; 
  signal FC1_CNT_4_RSTF_PT_0 : STD_LOGIC; 
  signal FC1_CNT_4_D1 : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_0 : STD_LOGIC; 
  signal EXP8_EXP : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_1 : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_2 : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_3 : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_4 : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_5 : STD_LOGIC; 
  signal FC1_CNT_4_D2 : STD_LOGIC; 
  signal FC1_CNT_4_D_TFF : STD_LOGIC; 
  signal FC1_CNT_5_EXP : STD_LOGIC; 
  signal EXP8_EXP_PT_0 : STD_LOGIC; 
  signal EXP8_EXP_PT_1 : STD_LOGIC; 
  signal EXP8_EXP_PT_2 : STD_LOGIC; 
  signal EXP8_EXP_PT_3 : STD_LOGIC; 
  signal EXP8_EXP_PT_4 : STD_LOGIC; 
  signal EXP8_EXP_PT_5 : STD_LOGIC; 
  signal FC1_CNT_5_Q : STD_LOGIC; 
  signal FC1_CNT_5_RSTF : STD_LOGIC; 
  signal FC1_CNT_5_R_OR_PRLD : STD_LOGIC; 
  signal FC1_CNT_5_D : STD_LOGIC; 
  signal FC1_CNT_5_RSTF_PT_0 : STD_LOGIC; 
  signal FC1_CNT_5_D1 : STD_LOGIC; 
  signal EXP7_EXP : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_0 : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_1 : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_2 : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_3 : STD_LOGIC; 
  signal FC1_CNT_5_D2 : STD_LOGIC; 
  signal FC1_CNT_5_D_TFF : STD_LOGIC; 
  signal FC1_CNT_5_EXP_PT_0 : STD_LOGIC; 
  signal EXP6_EXP : STD_LOGIC; 
  signal EXP7_EXP_PT_0 : STD_LOGIC; 
  signal EXP7_EXP_PT_1 : STD_LOGIC; 
  signal EXP7_EXP_PT_2 : STD_LOGIC; 
  signal EXP7_EXP_PT_3 : STD_LOGIC; 
  signal EXP7_EXP_PT_4 : STD_LOGIC; 
  signal EXP7_EXP_PT_5 : STD_LOGIC; 
  signal EXP6_EXP_PT_0 : STD_LOGIC; 
  signal EXP6_EXP_PT_1 : STD_LOGIC; 
  signal EXP6_EXP_PT_2 : STD_LOGIC; 
  signal EXP6_EXP_PT_3 : STD_LOGIC; 
  signal LIGHT_VALUE_3_Q : STD_LOGIC; 
  signal LIGHT_VALUE_3_D : STD_LOGIC; 
  signal LIGHT_VALUE_3_SETF : STD_LOGIC; 
  signal LIGHT_VALUE_3_SETF_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_3_D1 : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1 : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_2 : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2 : STD_LOGIC; 
  signal LIGHT_VALUE_3_D_TFF : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_1 : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP : STD_LOGIC; 
  signal FC1_CNT_6_Q : STD_LOGIC; 
  signal FC1_CNT_6_RSTF : STD_LOGIC; 
  signal FC1_CNT_6_R_OR_PRLD : STD_LOGIC; 
  signal FC1_CNT_6_D : STD_LOGIC; 
  signal FC1_CNT_6_RSTF_PT_0 : STD_LOGIC; 
  signal FC1_CNT_6_D1 : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_0 : STD_LOGIC; 
  signal EXP5_EXP : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_1 : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_2 : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_3 : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_4 : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_5 : STD_LOGIC; 
  signal FC1_CNT_6_D2 : STD_LOGIC; 
  signal FC1_CNT_6_D_TFF : STD_LOGIC; 
  signal EXP5_EXP_PT_0 : STD_LOGIC; 
  signal EXP5_EXP_PT_1 : STD_LOGIC; 
  signal EXP5_EXP_PT_2 : STD_LOGIC; 
  signal EXP5_EXP_PT_3 : STD_LOGIC; 
  signal EXP5_EXP_PT_4 : STD_LOGIC; 
  signal LIGHT_VALUE_0_Q : STD_LOGIC; 
  signal LIGHT_VALUE_0_RSTF : STD_LOGIC; 
  signal LIGHT_VALUE_0_R_OR_PRLD : STD_LOGIC; 
  signal LIGHT_VALUE_0_D : STD_LOGIC; 
  signal LIGHT_VALUE_0_RSTF_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_0_D1 : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_0 : STD_LOGIC; 
  signal TD1_CNT_5_EXP : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_1 : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_2 : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_3 : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_4 : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_5 : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2 : STD_LOGIC; 
  signal LIGHT_VALUE_0_D_TFF : STD_LOGIC; 
  signal TD1_CNT_5_Q : STD_LOGIC; 
  signal TD1_CNT_5_D : STD_LOGIC; 
  signal TD1_CNT_5_SETF : STD_LOGIC; 
  signal TD1_CNT_5_SETF_PT_0 : STD_LOGIC; 
  signal TD1_CNT_5_D1 : STD_LOGIC; 
  signal TD1_CNT_1_Q_3 : STD_LOGIC; 
  signal TD1_CNT_2_FBK : STD_LOGIC; 
  signal TD1_CNT_3_FBK : STD_LOGIC; 
  signal TD1_CNT_4_FBK : STD_LOGIC; 
  signal TD1_CNT_5_D2_PT_0 : STD_LOGIC; 
  signal TD1_CNT_5_D2 : STD_LOGIC; 
  signal TD1_CNT_5_D_TFF : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_0 : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_1 : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_2 : STD_LOGIC; 
  signal TD1_CNT_1_Q : STD_LOGIC; 
  signal TD1_CNT_1_D : STD_LOGIC; 
  signal TD1_CNT_1_SETF : STD_LOGIC; 
  signal TD1_CNT_1_SETF_PT_0 : STD_LOGIC; 
  signal TD1_CNT_1_D1 : STD_LOGIC; 
  signal TD1_CNT_1_D2_PT_0 : STD_LOGIC; 
  signal TD1_CNT_1_D2 : STD_LOGIC; 
  signal TD1_CNT_1_D_TFF : STD_LOGIC; 
  signal TD1_CNT_2_Q : STD_LOGIC; 
  signal TD1_CNT_2_RSTF : STD_LOGIC; 
  signal TD1_CNT_2_R_OR_PRLD : STD_LOGIC; 
  signal TD1_CNT_2_D : STD_LOGIC; 
  signal TD1_CNT_2_RSTF_PT_0 : STD_LOGIC; 
  signal TD1_CNT_2_D1 : STD_LOGIC; 
  signal TD1_CNT_2_D2_PT_0 : STD_LOGIC; 
  signal TD1_CNT_2_D2 : STD_LOGIC; 
  signal TD1_CNT_2_D_TFF : STD_LOGIC; 
  signal TD1_CNT_3_EXP_PT_0 : STD_LOGIC; 
  signal TD1_CNT_3_EXP_PT_1 : STD_LOGIC; 
  signal TD1_CNT_3_EXP : STD_LOGIC; 
  signal TD1_CNT_3_Q : STD_LOGIC; 
  signal TD1_CNT_3_D : STD_LOGIC; 
  signal TD1_CNT_3_SETF : STD_LOGIC; 
  signal TD1_CNT_3_SETF_PT_0 : STD_LOGIC; 
  signal TD1_CNT_3_D1 : STD_LOGIC; 
  signal TD1_CNT_3_D2_PT_0 : STD_LOGIC; 
  signal TD1_CNT_3_D2 : STD_LOGIC; 
  signal TD1_CNT_3_D_TFF : STD_LOGIC; 
  signal LIGHT_VALUE_2_Q : STD_LOGIC; 
  signal LIGHT_VALUE_2_RSTF : STD_LOGIC; 
  signal LIGHT_VALUE_2_R_OR_PRLD : STD_LOGIC; 
  signal LIGHT_VALUE_2_D : STD_LOGIC; 
  signal LIGHT_VALUE_2_RSTF_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_2_D1 : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_0 : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_1 : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_2 : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_3 : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_4 : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2 : STD_LOGIC; 
  signal LIGHT_VALUE_2_D_TFF : STD_LOGIC; 
  signal TD1_CNT_4_Q : STD_LOGIC; 
  signal TD1_CNT_4_RSTF : STD_LOGIC; 
  signal TD1_CNT_4_R_OR_PRLD : STD_LOGIC; 
  signal TD1_CNT_4_D : STD_LOGIC; 
  signal TD1_CNT_4_RSTF_PT_0 : STD_LOGIC; 
  signal TD1_CNT_4_D1 : STD_LOGIC; 
  signal TD1_CNT_4_D2_PT_0 : STD_LOGIC; 
  signal TD1_CNT_4_D2 : STD_LOGIC; 
  signal TD1_CNT_4_D_TFF : STD_LOGIC; 
  signal TD1_CNT_4_EXP_PT_0 : STD_LOGIC; 
  signal TD1_CNT_4_EXP_PT_1 : STD_LOGIC; 
  signal TD1_CNT_4_EXP_PT_2 : STD_LOGIC; 
  signal TD1_CNT_4_EXP : STD_LOGIC; 
  signal CM_FADE_UP_Q : STD_LOGIC; 
  signal CM_FADE_UP_R_OR_PRLD : STD_LOGIC; 
  signal CM_FADE_UP_D : STD_LOGIC; 
  signal CM_FADE_UP_D1 : STD_LOGIC; 
  signal CM_FADE_UP_D2_PT_0 : STD_LOGIC; 
  signal CM_FADE_UP_D2_PT_1 : STD_LOGIC; 
  signal CM_FADE_UP_D2_PT_2 : STD_LOGIC; 
  signal EXP15_EXP : STD_LOGIC; 
  signal CM_FADE_UP_D2_PT_3 : STD_LOGIC; 
  signal CM_FADE_UP_D2_PT_4 : STD_LOGIC; 
  signal CM_FADE_UP_D2_PT_5 : STD_LOGIC; 
  signal CM_FADE_UP_D2_PT_6 : STD_LOGIC; 
  signal CM_FADE_UP_D2 : STD_LOGIC; 
  signal CM_FADE_UP_D_TFF : STD_LOGIC; 
  signal CM_FADE_UP_FBK : STD_LOGIC; 
  signal EXP16_EXP : STD_LOGIC; 
  signal EXP15_EXP_PT_0 : STD_LOGIC; 
  signal EXP15_EXP_PT_1 : STD_LOGIC; 
  signal EXP15_EXP_PT_2 : STD_LOGIC; 
  signal EXP15_EXP_PT_3 : STD_LOGIC; 
  signal EXP15_EXP_PT_4 : STD_LOGIC; 
  signal EXP15_EXP_PT_5 : STD_LOGIC; 
  signal EXP16_EXP_PT_0 : STD_LOGIC; 
  signal EXP16_EXP_PT_1 : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_Q : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D1 : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_0 : STD_LOGIC; 
  signal EXP11_EXP : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_1 : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_2 : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_3 : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_4 : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_5 : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_6 : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2 : STD_LOGIC; 
  signal EXP11_EXP_PT_0 : STD_LOGIC; 
  signal EXP11_EXP_PT_1 : STD_LOGIC; 
  signal EXP11_EXP_PT_2 : STD_LOGIC; 
  signal EXP11_EXP_PT_3 : STD_LOGIC; 
  signal EXP11_EXP_PT_4 : STD_LOGIC; 
  signal EXP11_EXP_PT_5 : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D2_PT_1_0_INV : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D2_PT_2_0_INV : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D2_PT_2_1_INV : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D2_PT_3_0_INV : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_D2_PT_4_0_INV : STD_LOGIC; 
  signal TD1_TRIAC_TRIG_I_XOR_0_INV : STD_LOGIC; 
  signal EXP1_EXP_PT_0_0_INV : STD_LOGIC; 
  signal EXP1_EXP_PT_0_1_INV : STD_LOGIC; 
  signal EXP1_EXP_PT_1_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_D2_PT_1_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_D2_PT_1_12_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_0_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_0_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_0_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_0_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_0_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_1_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_1_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_1_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_1_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_1_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_2_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_2_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_4_EXP_PT_2_7_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_0_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_2_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_3_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_4_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_5_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_6_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_7_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_8_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_9_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_10_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_11_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_13_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_0_14_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_1_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_2_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_3_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_4_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_5_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_6_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_7_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_9_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_10_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_11_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_13_INV : STD_LOGIC; 
  signal EXP0_EXP_PT_1_14_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_0_1_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_1_1_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_1_2_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_1_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_5_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_6_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_7_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_0_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_1_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_2_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_3_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_4_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_5_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_6_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_7_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_8_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_9_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_10_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_11_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_12_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_14_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_15_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_16_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_0_2_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_1_2_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_2_5_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_2_6_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_2_7_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_1_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_2_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_3_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_4_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_5_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_6_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_7_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_8_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_9_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_10_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_11_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_12_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_14_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_15_INV : STD_LOGIC; 
  signal EXP2_EXP_PT_3_16_INV : STD_LOGIC; 
  signal CM_FADE_DOWN_D2_PT_2_0_INV : STD_LOGIC; 
  signal CM_FADE_DOWN_D2_PT_2_1_INV : STD_LOGIC; 
  signal CM_FADE_DOWN_D2_PT_5_1_INV : STD_LOGIC; 
  signal CM_FADE_DOWN_D2_PT_6_0_INV : STD_LOGIC; 
  signal CM_FADE_DOWN_XOR_0_INV : STD_LOGIC; 
  signal RXD_READY_EXP_PT_0_1_INV : STD_LOGIC; 
  signal RXD_READY_EXP_PT_1_0_INV : STD_LOGIC; 
  signal RXD_READY_EXP_PT_2_1_INV : STD_LOGIC; 
  signal RXD_READY_EXP_PT_3_0_INV : STD_LOGIC; 
  signal RXD_READY_EXP_PT_4_1_INV : STD_LOGIC; 
  signal RXD_7_EXP_PT_0_1_INV : STD_LOGIC; 
  signal RXD_7_EXP_PT_1_0_INV : STD_LOGIC; 
  signal RXD_7_D2_PT_0_1_INV : STD_LOGIC; 
  signal RXD_7_D2_PT_0_3_INV : STD_LOGIC; 
  signal RXD_7_D2_PT_1_1_INV : STD_LOGIC; 
  signal RXD_7_D2_PT_1_2_INV : STD_LOGIC; 
  signal UAR1_BYTE_AVAIL_D2_PT_0_2_INV : STD_LOGIC; 
  signal UAR1_BYTE_AVAIL_D2_PT_0_3_INV : STD_LOGIC; 
  signal UAR1_BYTE_AVAIL_D2_PT_0_4_INV : STD_LOGIC; 
  signal UAR1_BIT_DONE_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BIT_DONE_D2_PT_0_1_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_2_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_2_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_2_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_2_4_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_2_5_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_2_6_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_3_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_3_1_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_3_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_3_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_3_5_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_3_6_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_4_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_4_1_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_4_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_4_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_4_5_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_4_6_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_5_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_5_1_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_5_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_5_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_5_5_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_5_6_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_6_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_6_1_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_6_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_6_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_6_5_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_D2_PT_6_6_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_11_XOR_0_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_0_1_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_0_5_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_1_1_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_1_2_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_1_3_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_1_4_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_1_5_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_2_4_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_2_5_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_3_1_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_3_2_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_3_3_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_3_4_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_3_6_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_4_1_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_4_2_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_4_3_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_4_4_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_4_5_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_4_6_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_4_7_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_4_8_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_4_9_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_4_10_INV : STD_LOGIC; 
  signal EXP9_EXP_PT_4_11_INV : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_0_D2_PT_1_0_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_3_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_3_D2_PT_0_1_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_3_D2_PT_1_0_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_0_1_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_0_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_1_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_2_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_0_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_1_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_3_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_4_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_XOR_0_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_1_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_1_D2_PT_0_1_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_2_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BM1_CURRENT_STATE_2_D2_PT_0_1_INV : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_1_D2_PT_1_0_INV : STD_LOGIC; 
  signal UAR1_BM1_SAMPLED_BITS_2_D2_PT_1_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_D2_PT_2_1_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_D2_PT_2_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_1_D2_PT_2_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_D2_PT_2_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_D2_PT_2_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_2_D2_PT_2_4_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_D2_PT_2_1_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_D2_PT_2_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_3_D2_PT_2_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_D2_PT_2_1_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_D2_PT_2_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_4_D2_PT_2_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_D2_PT_2_1_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_D2_PT_2_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_5_D2_PT_2_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_D2_PT_2_1_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_D2_PT_2_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_6_D2_PT_2_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_D2_PT_2_1_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_D2_PT_2_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_7_D2_PT_2_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_D2_PT_2_1_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_D2_PT_2_2_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_8_D2_PT_2_3_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_9_D2_PT_0_0_INV : STD_LOGIC; 
  signal UAR1_BC1_CURRENT_STATE_10_D2_PT_1_0_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_0_0_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_0_2_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_1_1_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_1_2_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_2_2_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_2_3_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_2_5_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_2_6_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_3_1_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_3_2_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_3_3_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_3_5_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_3_6_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_4_0_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_4_1_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_4_2_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_4_3_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_4_5_INV : STD_LOGIC; 
  signal EXP10_EXP_PT_4_6_INV : STD_LOGIC; 
  signal UAR1_BYTE_OUT_7_D2_PT_0_0_INV : STD_LOGIC; 
  signal RXD_5_D2_PT_0_1_INV : STD_LOGIC; 
  signal RXD_5_D2_PT_0_3_INV : STD_LOGIC; 
  signal RXD_5_D2_PT_1_1_INV : STD_LOGIC; 
  signal RXD_5_D2_PT_1_2_INV : STD_LOGIC; 
  signal UAR1_BYTE_OUT_5_D2_PT_0_0_INV : STD_LOGIC; 
  signal RXD_6_D2_PT_0_1_INV : STD_LOGIC; 
  signal RXD_6_D2_PT_0_3_INV : STD_LOGIC; 
  signal RXD_6_D2_PT_1_1_INV : STD_LOGIC; 
  signal RXD_6_D2_PT_1_2_INV : STD_LOGIC; 
  signal UAR1_BYTE_OUT_6_D2_PT_0_0_INV : STD_LOGIC; 
  signal RXD_2_D2_PT_0_1_INV : STD_LOGIC; 
  signal RXD_2_D2_PT_0_3_INV : STD_LOGIC; 
  signal RXD_2_D2_PT_1_1_INV : STD_LOGIC; 
  signal RXD_2_D2_PT_1_2_INV : STD_LOGIC; 
  signal UAR1_BYTE_OUT_2_D2_PT_0_0_INV : STD_LOGIC; 
  signal EXP19_EXP_PT_0_1_INV : STD_LOGIC; 
  signal EXP19_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP19_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP19_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP19_EXP_PT_4_1_INV : STD_LOGIC; 
  signal EXP20_EXP_PT_1_1_INV : STD_LOGIC; 
  signal EXP20_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP20_EXP_PT_4_0_INV : STD_LOGIC; 
  signal EXP20_EXP_PT_4_1_INV : STD_LOGIC; 
  signal EXP20_EXP_PT_5_0_INV : STD_LOGIC; 
  signal RXD_1_EXP_PT_1_0_INV : STD_LOGIC; 
  signal RXD_1_EXP_PT_1_2_INV : STD_LOGIC; 
  signal RXD_1_D2_PT_0_1_INV : STD_LOGIC; 
  signal RXD_1_D2_PT_0_3_INV : STD_LOGIC; 
  signal RXD_1_D2_PT_1_1_INV : STD_LOGIC; 
  signal RXD_1_D2_PT_1_2_INV : STD_LOGIC; 
  signal UAR1_BYTE_OUT_1_D2_PT_0_0_INV : STD_LOGIC; 
  signal RXD_3_D2_PT_0_2_INV : STD_LOGIC; 
  signal RXD_3_D2_PT_0_3_INV : STD_LOGIC; 
  signal RXD_3_D2_PT_1_0_INV : STD_LOGIC; 
  signal RXD_3_D2_PT_1_2_INV : STD_LOGIC; 
  signal UAR1_BYTE_OUT_3_D2_PT_0_0_INV : STD_LOGIC; 
  signal RXD_0_EXP_PT_1_0_INV : STD_LOGIC; 
  signal RXD_0_EXP_PT_1_2_INV : STD_LOGIC; 
  signal RXD_0_D2_PT_0_1_INV : STD_LOGIC; 
  signal RXD_0_D2_PT_0_3_INV : STD_LOGIC; 
  signal RXD_0_D2_PT_1_1_INV : STD_LOGIC; 
  signal RXD_0_D2_PT_1_2_INV : STD_LOGIC; 
  signal UAR1_BYTE_OUT_0_D2_PT_0_0_INV : STD_LOGIC; 
  signal CM_PANIC_ON_D2_PT_4_0_INV : STD_LOGIC; 
  signal CM_PANIC_ON_D2_PT_4_1_INV : STD_LOGIC; 
  signal CM_PANIC_ON_D2_PT_5_1_INV : STD_LOGIC; 
  signal CM_PANIC_ON_D2_PT_6_0_INV : STD_LOGIC; 
  signal CM_PANIC_ON_XOR_0_INV : STD_LOGIC; 
  signal EXP17_EXP_PT_0_1_INV : STD_LOGIC; 
  signal EXP17_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP17_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP17_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP17_EXP_PT_4_1_INV : STD_LOGIC; 
  signal EXP18_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP18_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP18_EXP_PT_3_1_INV : STD_LOGIC; 
  signal EXP18_EXP_PT_4_0_INV : STD_LOGIC; 
  signal EXP18_EXP_PT_5_0_INV : STD_LOGIC; 
  signal RXD_4_D2_PT_0_1_INV : STD_LOGIC; 
  signal RXD_4_D2_PT_0_3_INV : STD_LOGIC; 
  signal RXD_4_D2_PT_1_1_INV : STD_LOGIC; 
  signal RXD_4_D2_PT_1_2_INV : STD_LOGIC; 
  signal UAR1_BYTE_OUT_4_D2_PT_0_0_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_1_0_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_1_1_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_XOR_0_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_0_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_2_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_3_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_4_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_5_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_6_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_7_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_8_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_0_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_1_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_2_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_3_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_4_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_5_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_6_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_7_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_1_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_9_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_10_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_1_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_9_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_10_INV : STD_LOGIC; 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_11_INV : STD_LOGIC; 
  signal FC1_CNT_3_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal FC1_CNT_3_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2_0_INV : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2_1_INV : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2_2_INV : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2_3_INV : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2_4_INV : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2_5_INV : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2_6_INV : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2_7_INV : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2_8_INV : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2_9_INV : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2_10_INV : STD_LOGIC; 
  signal FC1_CNT_3_D2_PT_2_11_INV : STD_LOGIC; 
  signal FC1_CNT_3_XOR_0_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_0_0_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_0_2_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_0_3_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_0_4_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_0_5_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_0_6_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_1_0_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_1_1_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_1_2_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_1_3_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_1_4_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_1_5_INV : STD_LOGIC; 
  signal FC1_CNT_3_EXP_PT_1_6_INV : STD_LOGIC; 
  signal EXP4_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP4_EXP_PT_3_1_INV : STD_LOGIC; 
  signal FC1_CNT_7_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal FC1_CNT_7_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_7_D2_PT_1_8_INV : STD_LOGIC; 
  signal FC1_CNT_7_D2_PT_1_9_INV : STD_LOGIC; 
  signal FC1_CNT_7_EXP_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_7_EXP_PT_1_0_INV : STD_LOGIC; 
  signal FC1_CNT_7_EXP_PT_1_1_INV : STD_LOGIC; 
  signal FC1_CNT_7_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_1_1_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_1_2_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_1_3_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_1_4_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_1_5_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_1_6_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_1_7_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_2_2_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_2_3_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_2_4_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_2_5_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_2_6_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_2_7_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_3_1_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_3_2_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_3_3_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_3_4_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_3_5_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_3_6_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_3_7_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_4_0_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_4_1_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_4_2_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_4_3_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_4_4_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_4_5_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_4_6_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_4_7_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_5_0_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_5_1_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_5_2_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_5_3_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_5_4_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_5_5_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_5_6_INV : STD_LOGIC; 
  signal EXP3_EXP_PT_5_7_INV : STD_LOGIC; 
  signal FC1_CNT_1_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal FC1_CNT_1_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_0_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_1_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_2_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_3_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_4_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_5_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_6_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_7_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_8_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_9_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_10_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_11_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_12_INV : STD_LOGIC; 
  signal FC1_CNT_1_D2_PT_4_13_INV : STD_LOGIC; 
  signal FC1_CNT_1_XOR_0_INV : STD_LOGIC; 
  signal FC1_CNT_0_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal FC1_CNT_0_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_0_XOR_0_INV : STD_LOGIC; 
  signal FC1_CNT_0_EXP_PT_1_0_INV : STD_LOGIC; 
  signal FC1_CNT_0_EXP_PT_1_1_INV : STD_LOGIC; 
  signal FC1_CNT_0_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_0_0_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_0_1_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_1_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_2_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_3_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_4_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_5_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_6_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_7_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_8_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_9_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_10_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_11_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_12_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_13_INV : STD_LOGIC; 
  signal EXP12_EXP_PT_4_14_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_SETF_PT_0_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_SETF_PT_0_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_D2_PT_1_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_D2_PT_1_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0_7_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0_10_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0_11_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0_12_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_0_13_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1_7_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1_10_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1_11_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_1_12_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_2_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_2_13_INV : STD_LOGIC; 
  signal LIGHT_VALUE_5_EXP_PT_2_14_INV : STD_LOGIC; 
  signal TD1_CNT_0_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_0_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_0_D2_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_0_D2_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_3_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_4_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_5_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_6_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_7_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_8_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_9_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_10_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_11_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_12_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_13_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_14_INV : STD_LOGIC; 
  signal TD1_CNT_0_EXP_PT_0_15_INV : STD_LOGIC; 
  signal TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_2_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal FC1_CNT_2_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_0_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_1_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_2_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_3_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_4_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_5_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_6_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_7_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_8_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_9_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_10_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_11_INV : STD_LOGIC; 
  signal FC1_CNT_2_D2_PT_2_12_INV : STD_LOGIC; 
  signal FC1_CNT_2_XOR_0_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_0_2_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_0_3_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_0_4_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_0_5_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_0_6_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_0_7_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_0_8_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_0_9_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_1_1_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_1_2_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_1_3_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_1_4_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_1_5_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_1_6_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_1_7_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_1_8_INV : STD_LOGIC; 
  signal FC1_CNT_2_EXP_PT_1_9_INV : STD_LOGIC; 
  signal EXP14_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP14_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP14_EXP_PT_3_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_SETF_PT_0_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_SETF_PT_0_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_1_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_1_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_1_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_1_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_1_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_1_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_1_7_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_1_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_1_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_1_11_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_2_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_2_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_2_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_2_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_2_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_2_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_2_7_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_2_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_2_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_2_11_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_3_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_D2_PT_3_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_1_EXP_PT_0_1_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_0_1_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_0_3_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_0_4_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_0_5_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_0_6_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_0_7_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_0_8_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_0_9_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_0_10_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_0_11_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_1_1_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_1_2_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_1_3_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_1_4_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_1_5_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_1_6_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_1_7_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_1_8_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_1_9_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_1_10_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_2_2_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_2_3_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_2_4_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_2_5_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_2_6_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_2_7_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_2_8_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_2_9_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_2_10_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_3_11_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_3_12_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_4_0_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_4_10_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_4_11_INV : STD_LOGIC; 
  signal EXP13_EXP_PT_4_13_INV : STD_LOGIC; 
  signal FC1_CNT_4_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal FC1_CNT_4_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_2_5_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_2_6_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_3_0_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_3_1_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_3_2_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_3_3_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_3_5_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_4_0_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_4_1_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_4_2_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_4_3_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_4_5_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_5_0_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_5_1_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_5_2_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_5_3_INV : STD_LOGIC; 
  signal FC1_CNT_4_D2_PT_5_4_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_1_1_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_1_2_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_1_3_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_1_5_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_2_2_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_2_3_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_2_4_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_3_1_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_3_2_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_3_3_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_3_4_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_4_0_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_4_1_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_4_2_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_4_3_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_4_4_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_5_0_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_5_1_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_5_2_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_5_3_INV : STD_LOGIC; 
  signal EXP8_EXP_PT_5_4_INV : STD_LOGIC; 
  signal FC1_CNT_5_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal FC1_CNT_5_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_1_6_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_1_7_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_2_0_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_2_1_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_2_2_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_2_3_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_2_4_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_2_6_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_3_0_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_3_1_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_3_2_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_3_3_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_3_4_INV : STD_LOGIC; 
  signal FC1_CNT_5_D2_PT_3_5_INV : STD_LOGIC; 
  signal FC1_CNT_5_EXP_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_5_EXP_PT_0_6_INV : STD_LOGIC; 
  signal FC1_CNT_5_EXP_PT_0_7_INV : STD_LOGIC; 
  signal FC1_CNT_5_EXP_PT_0_8_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_1_1_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_1_2_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_1_3_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_1_4_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_1_6_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_2_2_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_2_3_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_2_4_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_2_5_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_3_1_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_3_2_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_3_3_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_3_4_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_3_5_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_4_0_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_4_1_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_4_2_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_4_3_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_4_4_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_4_5_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_5_0_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_5_1_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_5_2_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_5_3_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_5_4_INV : STD_LOGIC; 
  signal EXP7_EXP_PT_5_5_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_0_0_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_0_2_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_0_3_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_0_4_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_0_5_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_0_6_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_1_1_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_1_2_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_1_3_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_1_4_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_1_5_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_2_7_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_2_8_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_3_1_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_3_7_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_3_8_INV : STD_LOGIC; 
  signal EXP6_EXP_PT_3_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_SETF_PT_0_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_SETF_PT_0_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1_7_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1_10_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1_11_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_1_12_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_2_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_D2_PT_2_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_0_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_0_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_0_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_0_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_0_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_0_7_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_0_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_0_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_0_10_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_0_11_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_0_12_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_1_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_1_12_INV : STD_LOGIC; 
  signal LIGHT_VALUE_3_EXP_PT_1_13_INV : STD_LOGIC; 
  signal FC1_CNT_6_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal FC1_CNT_6_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_2_7_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_2_8_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_3_0_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_3_1_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_3_2_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_3_3_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_3_4_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_3_5_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_3_7_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_4_0_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_4_1_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_4_2_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_4_3_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_4_4_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_4_5_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_4_6_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_5_0_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_5_1_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_5_2_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_5_3_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_5_4_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_5_5_INV : STD_LOGIC; 
  signal FC1_CNT_6_D2_PT_5_6_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_0_0_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_0_2_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_0_3_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_0_4_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_0_5_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_0_6_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_0_7_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_1_1_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_1_2_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_1_3_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_1_4_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_1_5_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_1_6_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_2_2_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_2_3_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_2_4_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_2_5_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_2_6_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_3_1_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_3_8_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_3_9_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_4_1_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_4_8_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_4_9_INV : STD_LOGIC; 
  signal EXP5_EXP_PT_4_10_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_2_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_2_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_2_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_2_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_2_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_2_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_2_7_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_2_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_2_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_3_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_3_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_3_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_3_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_3_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_3_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_3_7_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_3_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_3_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_4_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_4_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_4_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_4_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_4_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_4_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_4_7_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_4_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_4_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_5_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_0_D2_PT_5_2_INV : STD_LOGIC; 
  signal TD1_CNT_5_SETF_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_5_SETF_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_5_D2_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_5_D2_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_5_D2_PT_0_2_INV : STD_LOGIC; 
  signal TD1_CNT_5_D2_PT_0_3_INV : STD_LOGIC; 
  signal TD1_CNT_5_D2_PT_0_4_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_0_3_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_0_4_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_0_5_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_0_6_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_0_7_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_0_8_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_0_9_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_0_10_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_1_0_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_1_10_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_1_11_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_2_0_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_2_10_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_2_11_INV : STD_LOGIC; 
  signal TD1_CNT_5_EXP_PT_2_12_INV : STD_LOGIC; 
  signal TD1_CNT_1_SETF_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_1_SETF_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_1_XOR_0_INV : STD_LOGIC; 
  signal TD1_CNT_2_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_2_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_2_D2_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_2_D2_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_3_EXP_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_3_EXP_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_3_EXP_PT_0_2_INV : STD_LOGIC; 
  signal TD1_CNT_3_EXP_PT_0_3_INV : STD_LOGIC; 
  signal TD1_CNT_3_EXP_PT_1_0_INV : STD_LOGIC; 
  signal TD1_CNT_3_EXP_PT_1_1_INV : STD_LOGIC; 
  signal TD1_CNT_3_EXP_PT_1_2_INV : STD_LOGIC; 
  signal TD1_CNT_3_SETF_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_3_SETF_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_3_D2_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_3_D2_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_3_D2_PT_0_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_1_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_1_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_1_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_1_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_1_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_1_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_1_7_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_1_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_1_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_1_10_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_1_12_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_2_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_2_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_2_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_2_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_2_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_2_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_2_7_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_2_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_2_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_2_10_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_2_11_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_3_1_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_3_2_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_3_3_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_3_4_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_3_5_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_3_6_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_3_7_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_3_8_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_3_9_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_3_10_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_3_11_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_4_0_INV : STD_LOGIC; 
  signal LIGHT_VALUE_2_D2_PT_4_2_INV : STD_LOGIC; 
  signal TD1_CNT_4_RSTF_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_4_RSTF_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_4_D2_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_4_D2_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_4_D2_PT_0_2_INV : STD_LOGIC; 
  signal TD1_CNT_4_D2_PT_0_3_INV : STD_LOGIC; 
  signal TD1_CNT_4_EXP_PT_0_0_INV : STD_LOGIC; 
  signal TD1_CNT_4_EXP_PT_0_1_INV : STD_LOGIC; 
  signal TD1_CNT_4_EXP_PT_0_2_INV : STD_LOGIC; 
  signal TD1_CNT_4_EXP_PT_1_0_INV : STD_LOGIC; 
  signal TD1_CNT_4_EXP_PT_1_1_INV : STD_LOGIC; 
  signal TD1_CNT_4_EXP_PT_2_0_INV : STD_LOGIC; 
  signal CM_FADE_UP_D2_PT_2_0_INV : STD_LOGIC; 
  signal CM_FADE_UP_D2_PT_2_1_INV : STD_LOGIC; 
  signal CM_FADE_UP_D2_PT_5_1_INV : STD_LOGIC; 
  signal CM_FADE_UP_D2_PT_6_0_INV : STD_LOGIC; 
  signal CM_FADE_UP_XOR_0_INV : STD_LOGIC; 
  signal EXP15_EXP_PT_1_1_INV : STD_LOGIC; 
  signal EXP15_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP15_EXP_PT_3_1_INV : STD_LOGIC; 
  signal EXP15_EXP_PT_4_1_INV : STD_LOGIC; 
  signal EXP15_EXP_PT_5_0_INV : STD_LOGIC; 
  signal EXP16_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP16_EXP_PT_1_1_INV : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_2_0_INV : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_3_0_INV : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_3_1_INV : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_4_0_INV : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_5_0_INV : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_5_1_INV : STD_LOGIC; 
  signal Q_OPTX_FX_DC_68_D2_PT_6_0_INV : STD_LOGIC; 
  signal EXP11_EXP_PT_1_0_INV : STD_LOGIC; 
  signal EXP11_EXP_PT_1_1_INV : STD_LOGIC; 
  signal EXP11_EXP_PT_1_2_INV : STD_LOGIC; 
  signal EXP11_EXP_PT_2_0_INV : STD_LOGIC; 
  signal EXP11_EXP_PT_2_1_INV : STD_LOGIC; 
  signal EXP11_EXP_PT_2_2_INV : STD_LOGIC; 
  signal EXP11_EXP_PT_3_0_INV : STD_LOGIC; 
  signal EXP11_EXP_PT_3_1_INV : STD_LOGIC; 
  signal EXP11_EXP_PT_4_0_INV : STD_LOGIC; 
  signal EXP11_EXP_PT_4_1_INV : STD_LOGIC; 
  signal EXP11_EXP_PT_5_0_INV : STD_LOGIC; 
  signal EXP11_EXP_PT_5_1_INV : STD_LOGIC; 
  signal GND : STD_LOGIC; 
  signal PRLD : STD_LOGIC; 
  signal VCC : STD_LOGIC; 
  signal LIGHT_VALUE : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal FC1_CNT : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal DFSM1_CURRENT_STATE_H_CURRENT_STATE : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal RC_ADDRESS_C : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal UAR1_BYTE_OUT : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal UAR1_BM1_SAMPLED_BITS : STD_LOGIC_VECTOR ( 2 downto 0 ); 
begin
  TRIAC_PULSE_9 : X_BUF 
    port map (
      I => TD1_TRIAC_TRIG_I,
      O => TRIAC_PULSE
    );
  TD1_TRIAC_TRIG_I_10 : X_BUF 
    port map (
      I => TD1_TRIAC_TRIG_I_Q,
      O => TD1_TRIAC_TRIG_I
    );
  TD1_TRIAC_TRIG_I_REG : X_BUF 
    port map (
      I => TD1_TRIAC_TRIG_I_D,
      O => TD1_TRIAC_TRIG_I_Q
    );
  GND_ZERO : X_ZERO 
    port map (
      O => GND
    );
  TD1_TRIAC_TRIG_I_D1_11 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => TD1_TRIAC_TRIG_I_D1
    );
  TD1_TRIAC_TRIG_I_D2_PT_0_12 : X_AND2 
    port map (
      I0 => EXP1_EXP,
      I1 => EXP1_EXP,
      O => TD1_TRIAC_TRIG_I_D2_PT_0
    );
  TD1_TRIAC_TRIG_I_D2_PT_1_13 : X_AND2 
    port map (
      I0 => TD1_TRIAC_TRIG_I_D2_PT_1_0_INV,
      I1 => TD1_CNT_5_Q_0,
      O => TD1_TRIAC_TRIG_I_D2_PT_1
    );
  TD1_TRIAC_TRIG_I_D2_PT_2_14 : X_AND3 
    port map (
      I0 => TD1_TRIAC_TRIG_I_D2_PT_2_0_INV,
      I1 => TD1_TRIAC_TRIG_I_D2_PT_2_1_INV,
      I2 => TD1_CNT_4_Q_1,
      O => TD1_TRIAC_TRIG_I_D2_PT_2
    );
  TD1_TRIAC_TRIG_I_D2_PT_3_15 : X_AND3 
    port map (
      I0 => TD1_TRIAC_TRIG_I_D2_PT_3_0_INV,
      I1 => TD1_CNT_4_Q_1,
      I2 => TD1_CNT_5_Q_0,
      O => TD1_TRIAC_TRIG_I_D2_PT_3
    );
  TD1_TRIAC_TRIG_I_D2_PT_4_16 : X_AND3 
    port map (
      I0 => TD1_TRIAC_TRIG_I_D2_PT_4_0_INV,
      I1 => TD1_CNT_5_Q_0,
      I2 => Q_OPTX_FX_DC_68_UIM,
      O => TD1_TRIAC_TRIG_I_D2_PT_4
    );
  TD1_TRIAC_TRIG_I_D2_PT_5_17 : X_AND3 
    port map (
      I0 => TD1_CNT_4_Q_1,
      I1 => TD1_CNT_5_Q_0,
      I2 => Q_OPTX_FX_DC_68_UIM,
      O => TD1_TRIAC_TRIG_I_D2_PT_5
    );
  TD1_TRIAC_TRIG_I_D2_18 : X_OR6 
    port map (
      I0 => TD1_TRIAC_TRIG_I_D2_PT_0,
      I1 => TD1_TRIAC_TRIG_I_D2_PT_1,
      I2 => TD1_TRIAC_TRIG_I_D2_PT_2,
      I3 => TD1_TRIAC_TRIG_I_D2_PT_3,
      I4 => TD1_TRIAC_TRIG_I_D2_PT_4,
      I5 => TD1_TRIAC_TRIG_I_D2_PT_5,
      O => TD1_TRIAC_TRIG_I_D2
    );
  TD1_TRIAC_TRIG_I_XOR : X_XOR2 
    port map (
      I0 => TD1_TRIAC_TRIG_I_XOR_0_INV,
      I1 => TD1_TRIAC_TRIG_I_D2,
      O => TD1_TRIAC_TRIG_I_D
    );
  EXP1_EXP_PT_0_19 : X_AND3 
    port map (
      I0 => EXP1_EXP_PT_0_0_INV,
      I1 => EXP1_EXP_PT_0_1_INV,
      I2 => Q_OPTX_FX_DC_68_UIM,
      O => EXP1_EXP_PT_0
    );
  EXP1_EXP_PT_1_20 : X_AND3 
    port map (
      I0 => EXP1_EXP_PT_1_0_INV,
      I1 => TD1_CNT_4_Q_1,
      I2 => Q_OPTX_FX_DC_68_UIM,
      O => EXP1_EXP_PT_1
    );
  EXP1_EXP_21 : X_OR2 
    port map (
      I0 => EXP1_EXP_PT_0,
      I1 => EXP1_EXP_PT_1,
      O => EXP1_EXP
    );
  LIGHT_VALUE_4_Q_22 : X_BUF 
    port map (
      I => LIGHT_VALUE_4_Q,
      O => LIGHT_VALUE(4)
    );
  LIGHT_VALUE_4_R_OR_PRLD_23 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_4_RSTF,
      I1 => PRLD,
      O => LIGHT_VALUE_4_R_OR_PRLD
    );
  LIGHT_VALUE_4_REG : X_FF 
    port map (
      I => LIGHT_VALUE_4_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => LIGHT_VALUE_4_R_OR_PRLD,
      O => LIGHT_VALUE_4_Q
    );
  VCC_ONE : X_ONE 
    port map (
      O => VCC
    );
  LIGHT_VALUE_4_RSTF_PT_0_24 : X_AND2 
    port map (
      I0 => LIGHT_VALUE_4_RSTF_PT_0_0_INV,
      I1 => LIGHT_VALUE_4_RSTF_PT_0_1_INV,
      O => LIGHT_VALUE_4_RSTF_PT_0
    );
  LIGHT_VALUE_4_RSTF_25 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_4_RSTF_PT_0,
      I1 => LIGHT_VALUE_4_RSTF_PT_0,
      O => LIGHT_VALUE_4_RSTF
    );
  LIGHT_VALUE_4_D1_26 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => LIGHT_VALUE_4_D1
    );
  LIGHT_VALUE_4_D2_PT_0_27 : X_AND2 
    port map (
      I0 => EXP0_EXP,
      I1 => EXP0_EXP,
      O => LIGHT_VALUE_4_D2_PT_0
    );
  LIGHT_VALUE_4_D2_PT_1_28 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => FC1_CNT_3_FBK,
      I2 => FC1_CNT(1),
      I3 => FC1_CNT(2),
      I4 => FC1_CNT_4_FBK,
      I5 => FC1_CNT_5_FBK,
      I6 => FC1_CNT_6_FBK,
      I7 => FC1_CNT(0),
      I8 => LIGHT_VALUE_4_D2_PT_1_8_INV,
      I9 => LIGHT_VALUE(3),
      I10 => LIGHT_VALUE(1),
      I11 => LIGHT_VALUE(2),
      I12 => LIGHT_VALUE_4_D2_PT_1_12_INV,
      I13 => LIGHT_VALUE(0),
      I14 => FC1_CNT_7_FBK,
      I15 => VCC,
      O => LIGHT_VALUE_4_D2_PT_1
    );
  LIGHT_VALUE_4_D2_29 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_4_D2_PT_0,
      I1 => LIGHT_VALUE_4_D2_PT_1,
      O => LIGHT_VALUE_4_D2
    );
  LIGHT_VALUE_4_D_30 : X_XOR2 
    port map (
      I0 => LIGHT_VALUE_4_D_TFF,
      I1 => LIGHT_VALUE_4_Q,
      O => LIGHT_VALUE_4_D
    );
  LIGHT_VALUE_4_XOR : X_XOR2 
    port map (
      I0 => LIGHT_VALUE_4_D1,
      I1 => LIGHT_VALUE_4_D2,
      O => LIGHT_VALUE_4_D_TFF
    );
  LIGHT_VALUE_4_EXP_PT_0_31 : X_AND7 
    port map (
      I0 => LIGHT_VALUE_4_EXP_PT_0_0_INV,
      I1 => LIGHT_VALUE_4_FBK,
      I2 => LIGHT_VALUE_4_EXP_PT_0_2_INV,
      I3 => LIGHT_VALUE_4_EXP_PT_0_3_INV,
      I4 => LIGHT_VALUE_4_EXP_PT_0_4_INV,
      I5 => LIGHT_VALUE_4_EXP_PT_0_5_INV,
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => LIGHT_VALUE_4_EXP_PT_0
    );
  LIGHT_VALUE_4_EXP_PT_1_32 : X_AND7 
    port map (
      I0 => LIGHT_VALUE_4_EXP_PT_1_0_INV,
      I1 => LIGHT_VALUE_4_EXP_PT_1_1_INV,
      I2 => LIGHT_VALUE_4_EXP_PT_1_2_INV,
      I3 => LIGHT_VALUE_4_EXP_PT_1_3_INV,
      I4 => LIGHT_VALUE_4_EXP_PT_1_4_INV,
      I5 => LIGHT_VALUE(5),
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => LIGHT_VALUE_4_EXP_PT_1
    );
  LIGHT_VALUE_4_EXP_PT_2_33 : X_AND8 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => LIGHT_VALUE_4_EXP_PT_2_1_INV,
      I2 => FC1_CNT_3_FBK,
      I3 => FC1_CNT(1),
      I4 => FC1_CNT(2),
      I5 => FC1_CNT(0),
      I6 => LIGHT_VALUE_4_EXP_PT_2_6_INV,
      I7 => LIGHT_VALUE_4_EXP_PT_2_7_INV,
      O => LIGHT_VALUE_4_EXP_PT_2
    );
  LIGHT_VALUE_4_EXP_34 : X_OR3 
    port map (
      I0 => LIGHT_VALUE_4_EXP_PT_0,
      I1 => LIGHT_VALUE_4_EXP_PT_1,
      I2 => LIGHT_VALUE_4_EXP_PT_2,
      O => LIGHT_VALUE_4_EXP
    );
  LIGHT_VALUE_4_FBK_35 : X_BUF 
    port map (
      I => LIGHT_VALUE_4_Q,
      O => LIGHT_VALUE_4_FBK
    );
  EXP0_EXP_PT_0_36 : X_AND16 
    port map (
      I0 => EXP0_EXP_PT_0_0_INV,
      I1 => LIGHT_VALUE_4_FBK,
      I2 => EXP0_EXP_PT_0_2_INV,
      I3 => EXP0_EXP_PT_0_3_INV,
      I4 => EXP0_EXP_PT_0_4_INV,
      I5 => EXP0_EXP_PT_0_5_INV,
      I6 => EXP0_EXP_PT_0_6_INV,
      I7 => EXP0_EXP_PT_0_7_INV,
      I8 => EXP0_EXP_PT_0_8_INV,
      I9 => EXP0_EXP_PT_0_9_INV,
      I10 => EXP0_EXP_PT_0_10_INV,
      I11 => EXP0_EXP_PT_0_11_INV,
      I12 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I13 => EXP0_EXP_PT_0_13_INV,
      I14 => EXP0_EXP_PT_0_14_INV,
      I15 => VCC,
      O => EXP0_EXP_PT_0
    );
  EXP0_EXP_PT_1_37 : X_AND16 
    port map (
      I0 => EXP0_EXP_PT_1_0_INV,
      I1 => EXP0_EXP_PT_1_1_INV,
      I2 => EXP0_EXP_PT_1_2_INV,
      I3 => EXP0_EXP_PT_1_3_INV,
      I4 => EXP0_EXP_PT_1_4_INV,
      I5 => EXP0_EXP_PT_1_5_INV,
      I6 => EXP0_EXP_PT_1_6_INV,
      I7 => EXP0_EXP_PT_1_7_INV,
      I8 => LIGHT_VALUE(5),
      I9 => EXP0_EXP_PT_1_9_INV,
      I10 => EXP0_EXP_PT_1_10_INV,
      I11 => EXP0_EXP_PT_1_11_INV,
      I12 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I13 => EXP0_EXP_PT_1_13_INV,
      I14 => EXP0_EXP_PT_1_14_INV,
      I15 => VCC,
      O => EXP0_EXP_PT_1
    );
  EXP0_EXP_38 : X_OR2 
    port map (
      I0 => EXP0_EXP_PT_0,
      I1 => EXP0_EXP_PT_1,
      O => EXP0_EXP
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_Q_39 : X_BUF 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_Q,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1)
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_R_OR_PRLD_40 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_R_OR_PRLD
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_REG : X_FF 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_R_OR_PRLD,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_Q
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D1_41 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D1
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D2_PT_0_42 : X_AND2 
    port map (
      I0 => EXP2_EXP,
      I1 => EXP2_EXP,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D2_PT_0
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D2_PT_1_43 : X_AND2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => CM_PANIC_ON,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D2_PT_1
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D2_44 : X_OR2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D2_PT_0,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D2_PT_1,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D2
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D_45 : X_XOR2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D_TFF,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_Q,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_XOR : X_XOR2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D1,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D2,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_D_TFF
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_0_46 : X_AND3 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_0_1_INV,
      I2 => CM_PANIC_ON,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_0
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_1_47 : X_AND3 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_1_1_INV,
      I2 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_1_2_INV,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_1
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_48 : X_AND8 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_1_INV,
      I2 => LIGHT_VALUE(5),
      I3 => LIGHT_VALUE(3),
      I4 => LIGHT_VALUE(1),
      I5 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_5_INV,
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_6_INV,
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_7_INV,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_49 : X_AND32 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_1_INV,
      I2 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_2_INV,
      I3 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_3_INV,
      I4 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_4_INV,
      I5 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_5_INV,
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_6_INV,
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_7_INV,
      I8 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_8_INV,
      I9 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_9_INV,
      I10 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_10_INV,
      I11 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_11_INV,
      I12 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_12_INV,
      I13 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I14 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_14_INV,
      I15 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_15_INV,
      I16 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_16_INV,
      I17 => VCC,
      I18 => VCC,
      I19 => VCC,
      I20 => VCC,
      I21 => VCC,
      I22 => VCC,
      I23 => VCC,
      I24 => VCC,
      I25 => VCC,
      I26 => VCC,
      I27 => VCC,
      I28 => VCC,
      I29 => VCC,
      I30 => VCC,
      I31 => VCC,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_50 : X_OR4 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_0,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_1,
      I2 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2,
      I3 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK_51 : X_BUF 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_Q,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK
    );
  EXP2_EXP_PT_0_52 : X_AND3 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => CM_FADE_DOWN,
      I2 => EXP2_EXP_PT_0_2_INV,
      O => EXP2_EXP_PT_0
    );
  EXP2_EXP_PT_1_53 : X_AND4 
    port map (
      I0 => EXP2_EXP_PT_1_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I2 => EXP2_EXP_PT_1_2_INV,
      I3 => CM_FADE_UP,
      O => EXP2_EXP_PT_1
    );
  EXP2_EXP_PT_2_54 : X_AND8 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => EXP2_EXP_PT_2_1_INV,
      I2 => LIGHT_VALUE(5),
      I3 => LIGHT_VALUE(3),
      I4 => LIGHT_VALUE(1),
      I5 => EXP2_EXP_PT_2_5_INV,
      I6 => EXP2_EXP_PT_2_6_INV,
      I7 => EXP2_EXP_PT_2_7_INV,
      O => EXP2_EXP_PT_2
    );
  EXP2_EXP_PT_3_55 : X_AND32 
    port map (
      I0 => EXP2_EXP_PT_3_0_INV,
      I1 => EXP2_EXP_PT_3_1_INV,
      I2 => EXP2_EXP_PT_3_2_INV,
      I3 => EXP2_EXP_PT_3_3_INV,
      I4 => EXP2_EXP_PT_3_4_INV,
      I5 => EXP2_EXP_PT_3_5_INV,
      I6 => EXP2_EXP_PT_3_6_INV,
      I7 => EXP2_EXP_PT_3_7_INV,
      I8 => EXP2_EXP_PT_3_8_INV,
      I9 => EXP2_EXP_PT_3_9_INV,
      I10 => EXP2_EXP_PT_3_10_INV,
      I11 => EXP2_EXP_PT_3_11_INV,
      I12 => EXP2_EXP_PT_3_12_INV,
      I13 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I14 => EXP2_EXP_PT_3_14_INV,
      I15 => EXP2_EXP_PT_3_15_INV,
      I16 => EXP2_EXP_PT_3_16_INV,
      I17 => VCC,
      I18 => VCC,
      I19 => VCC,
      I20 => VCC,
      I21 => VCC,
      I22 => VCC,
      I23 => VCC,
      I24 => VCC,
      I25 => VCC,
      I26 => VCC,
      I27 => VCC,
      I28 => VCC,
      I29 => VCC,
      I30 => VCC,
      I31 => VCC,
      O => EXP2_EXP_PT_3
    );
  EXP2_EXP_56 : X_OR4 
    port map (
      I0 => EXP2_EXP_PT_0,
      I1 => EXP2_EXP_PT_1,
      I2 => EXP2_EXP_PT_2,
      I3 => EXP2_EXP_PT_3,
      O => EXP2_EXP
    );
  CM_FADE_DOWN_57 : X_BUF 
    port map (
      I => CM_FADE_DOWN_Q,
      O => CM_FADE_DOWN
    );
  CM_FADE_DOWN_R_OR_PRLD_58 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => CM_FADE_DOWN_R_OR_PRLD
    );
  CM_FADE_DOWN_REG : X_FF 
    port map (
      I => CM_FADE_DOWN_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => CM_FADE_DOWN_R_OR_PRLD,
      O => CM_FADE_DOWN_Q
    );
  CM_FADE_DOWN_D1_59 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => CM_FADE_DOWN_D1
    );
  CM_FADE_DOWN_D2_PT_0_60 : X_AND2 
    port map (
      I0 => RXD_ACK,
      I1 => RXD_ACK,
      O => CM_FADE_DOWN_D2_PT_0
    );
  CM_FADE_DOWN_D2_PT_1_61 : X_AND2 
    port map (
      I0 => RXD_2_FBK,
      I1 => RXD_2_FBK,
      O => CM_FADE_DOWN_D2_PT_1
    );
  CM_FADE_DOWN_D2_PT_2_62 : X_AND2 
    port map (
      I0 => CM_FADE_DOWN_D2_PT_2_0_INV,
      I1 => CM_FADE_DOWN_D2_PT_2_1_INV,
      O => CM_FADE_DOWN_D2_PT_2
    );
  CM_FADE_DOWN_D2_PT_3_63 : X_AND2 
    port map (
      I0 => EXP19_EXP,
      I1 => EXP19_EXP,
      O => CM_FADE_DOWN_D2_PT_3
    );
  CM_FADE_DOWN_D2_PT_4_64 : X_AND2 
    port map (
      I0 => EXP20_EXP,
      I1 => EXP20_EXP,
      O => CM_FADE_DOWN_D2_PT_4
    );
  CM_FADE_DOWN_D2_PT_5_65 : X_AND2 
    port map (
      I0 => RC_ADDRESS_C(0),
      I1 => CM_FADE_DOWN_D2_PT_5_1_INV,
      O => CM_FADE_DOWN_D2_PT_5
    );
  CM_FADE_DOWN_D2_PT_6_66 : X_AND2 
    port map (
      I0 => CM_FADE_DOWN_D2_PT_6_0_INV,
      I1 => RXD_4_FBK,
      O => CM_FADE_DOWN_D2_PT_6
    );
  CM_FADE_DOWN_D2_67 : X_OR7 
    port map (
      I0 => CM_FADE_DOWN_D2_PT_0,
      I1 => CM_FADE_DOWN_D2_PT_1,
      I2 => CM_FADE_DOWN_D2_PT_2,
      I3 => CM_FADE_DOWN_D2_PT_3,
      I4 => CM_FADE_DOWN_D2_PT_4,
      I5 => CM_FADE_DOWN_D2_PT_5,
      I6 => CM_FADE_DOWN_D2_PT_6,
      O => CM_FADE_DOWN_D2
    );
  CM_FADE_DOWN_D_68 : X_XOR2 
    port map (
      I0 => CM_FADE_DOWN_D_TFF,
      I1 => CM_FADE_DOWN_Q,
      O => CM_FADE_DOWN_D
    );
  CM_FADE_DOWN_XOR : X_XOR2 
    port map (
      I0 => CM_FADE_DOWN_XOR_0_INV,
      I1 => CM_FADE_DOWN_D2,
      O => CM_FADE_DOWN_D_TFF
    );
  CM_FADE_DOWN_FBK_69 : X_BUF 
    port map (
      I => CM_FADE_DOWN_Q,
      O => CM_FADE_DOWN_FBK
    );
  RXD_ACK_70 : X_BUF 
    port map (
      I => RXD_ACK_Q,
      O => RXD_ACK
    );
  RXD_ACK_R_OR_PRLD_71 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => RXD_ACK_R_OR_PRLD
    );
  RXD_ACK_REG : X_FF 
    port map (
      I => RXD_ACK_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => RXD_ACK_R_OR_PRLD,
      O => RXD_ACK_Q
    );
  RXD_ACK_D1_72 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => RXD_ACK_D1
    );
  RXD_ACK_D2_PT_0_73 : X_AND2 
    port map (
      I0 => RXD_READY,
      I1 => RXD_READY,
      O => RXD_ACK_D2_PT_0
    );
  RXD_ACK_D2_74 : X_OR2 
    port map (
      I0 => RXD_ACK_D2_PT_0,
      I1 => RXD_ACK_D2_PT_0,
      O => RXD_ACK_D2
    );
  RXD_ACK_XOR : X_XOR2 
    port map (
      I0 => RXD_ACK_D1,
      I1 => RXD_ACK_D2,
      O => RXD_ACK_D
    );
  RXD_READY_75 : X_BUF 
    port map (
      I => RXD_READY_Q,
      O => RXD_READY
    );
  RXD_READY_R_OR_PRLD_76 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => RXD_READY_R_OR_PRLD
    );
  RXD_READY_REG : X_FF 
    port map (
      I => RXD_READY_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => RXD_READY_R_OR_PRLD,
      O => RXD_READY_Q
    );
  RXD_READY_D1_77 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => RXD_READY_D1
    );
  RXD_READY_D2_PT_0_78 : X_AND2 
    port map (
      I0 => RXD_7_EXP,
      I1 => RXD_7_EXP,
      O => RXD_READY_D2_PT_0
    );
  RXD_READY_D2_79 : X_OR2 
    port map (
      I0 => RXD_READY_D2_PT_0,
      I1 => RXD_READY_D2_PT_0,
      O => RXD_READY_D2
    );
  RXD_READY_XOR : X_XOR2 
    port map (
      I0 => RXD_READY_D1,
      I1 => RXD_READY_D2,
      O => RXD_READY_D
    );
  RXD_READY_EXP_PT_0_80 : X_AND2 
    port map (
      I0 => RC_ADDRESS_C(1),
      I1 => RXD_READY_EXP_PT_0_1_INV,
      O => RXD_READY_EXP_PT_0
    );
  RXD_READY_EXP_PT_1_81 : X_AND2 
    port map (
      I0 => RXD_READY_EXP_PT_1_0_INV,
      I1 => RXD_5_FBK,
      O => RXD_READY_EXP_PT_1
    );
  RXD_READY_EXP_PT_2_82 : X_AND2 
    port map (
      I0 => RC_ADDRESS_C(2),
      I1 => RXD_READY_EXP_PT_2_1_INV,
      O => RXD_READY_EXP_PT_2
    );
  RXD_READY_EXP_PT_3_83 : X_AND2 
    port map (
      I0 => RXD_READY_EXP_PT_3_0_INV,
      I1 => RXD_6_FBK,
      O => RXD_READY_EXP_PT_3
    );
  RXD_READY_EXP_PT_4_84 : X_AND2 
    port map (
      I0 => RC_ADDRESS_C(3),
      I1 => RXD_READY_EXP_PT_4_1_INV,
      O => RXD_READY_EXP_PT_4
    );
  RXD_READY_EXP_85 : X_OR5 
    port map (
      I0 => RXD_READY_EXP_PT_0,
      I1 => RXD_READY_EXP_PT_1,
      I2 => RXD_READY_EXP_PT_2,
      I3 => RXD_READY_EXP_PT_3,
      I4 => RXD_READY_EXP_PT_4,
      O => RXD_READY_EXP
    );
  RXD_READY_FBK_86 : X_BUF 
    port map (
      I => RXD_READY_Q,
      O => RXD_READY_FBK
    );
  RXD_7_EXP_PT_0_87 : X_AND2 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_7_EXP_PT_0_1_INV,
      O => RXD_7_EXP_PT_0
    );
  RXD_7_EXP_PT_1_88 : X_AND2 
    port map (
      I0 => RXD_7_EXP_PT_1_0_INV,
      I1 => RXD_READY_FBK,
      O => RXD_7_EXP_PT_1
    );
  RXD_7_EXP_89 : X_OR2 
    port map (
      I0 => RXD_7_EXP_PT_0,
      I1 => RXD_7_EXP_PT_1,
      O => RXD_7_EXP
    );
  RXD_7_FBK_90 : X_BUF 
    port map (
      I => RXD_7_Q,
      O => RXD_7_FBK
    );
  RXD_7_R_OR_PRLD_91 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => RXD_7_R_OR_PRLD
    );
  RXD_7_REG : X_FF 
    port map (
      I => RXD_7_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => RXD_7_R_OR_PRLD,
      O => RXD_7_Q
    );
  RXD_7_D1_92 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => RXD_7_D1
    );
  RXD_7_D2_PT_0_93 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_7_D2_PT_0_1_INV,
      I2 => RXD_7_FBK,
      I3 => RXD_7_D2_PT_0_3_INV,
      O => RXD_7_D2_PT_0
    );
  RXD_7_D2_PT_1_94 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_7_D2_PT_1_1_INV,
      I2 => RXD_7_D2_PT_1_2_INV,
      I3 => UAR1_BYTE_OUT(7),
      O => RXD_7_D2_PT_1
    );
  RXD_7_D2_95 : X_OR2 
    port map (
      I0 => RXD_7_D2_PT_0,
      I1 => RXD_7_D2_PT_1,
      O => RXD_7_D2
    );
  RXD_7_D_96 : X_XOR2 
    port map (
      I0 => RXD_7_D_TFF,
      I1 => RXD_7_Q,
      O => RXD_7_D
    );
  RXD_7_XOR : X_XOR2 
    port map (
      I0 => RXD_7_D1,
      I1 => RXD_7_D2,
      O => RXD_7_D_TFF
    );
  UAR1_BYTE_AVAIL_97 : X_BUF 
    port map (
      I => UAR1_BYTE_AVAIL_Q,
      O => UAR1_BYTE_AVAIL
    );
  UAR1_BYTE_AVAIL_R_OR_PRLD_98 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BYTE_AVAIL_R_OR_PRLD
    );
  UAR1_BYTE_AVAIL_REG : X_FF 
    port map (
      I => UAR1_BYTE_AVAIL_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BYTE_AVAIL_R_OR_PRLD,
      O => UAR1_BYTE_AVAIL_Q
    );
  UAR1_BYTE_AVAIL_D1_99 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BYTE_AVAIL_D1
    );
  UAR1_BYTE_AVAIL_D2_PT_0_100 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE_FBK,
      I1 => UAR1_BC1_CURRENT_STATE_1_Q_4,
      I2 => UAR1_BYTE_AVAIL_D2_PT_0_2_INV,
      I3 => UAR1_BYTE_AVAIL_D2_PT_0_3_INV,
      I4 => UAR1_BYTE_AVAIL_D2_PT_0_4_INV,
      O => UAR1_BYTE_AVAIL_D2_PT_0
    );
  UAR1_BYTE_AVAIL_D2_101 : X_OR2 
    port map (
      I0 => UAR1_BYTE_AVAIL_D2_PT_0,
      I1 => UAR1_BYTE_AVAIL_D2_PT_0,
      O => UAR1_BYTE_AVAIL_D2
    );
  UAR1_BYTE_AVAIL_XOR : X_XOR2 
    port map (
      I0 => UAR1_BYTE_AVAIL_D1,
      I1 => UAR1_BYTE_AVAIL_D2,
      O => UAR1_BYTE_AVAIL_D
    );
  UAR1_BYTE_AVAIL_FBK_102 : X_BUF 
    port map (
      I => UAR1_BYTE_AVAIL_Q,
      O => UAR1_BYTE_AVAIL_FBK
    );
  UAR1_BIT_DONE_103 : X_BUF 
    port map (
      I => UAR1_BIT_DONE_Q,
      O => UAR1_BIT_DONE
    );
  UAR1_BIT_DONE_R_OR_PRLD_104 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BIT_DONE_R_OR_PRLD
    );
  UAR1_BIT_DONE_REG : X_FF 
    port map (
      I => UAR1_BIT_DONE_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BIT_DONE_R_OR_PRLD,
      O => UAR1_BIT_DONE_Q
    );
  UAR1_BIT_DONE_D1_105 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BIT_DONE_D1
    );
  UAR1_BIT_DONE_D2_PT_0_106 : X_AND3 
    port map (
      I0 => UAR1_BIT_DONE_D2_PT_0_0_INV,
      I1 => UAR1_BIT_DONE_D2_PT_0_1_INV,
      I2 => UAR1_BM1_CURRENT_STATE_1_FBK,
      O => UAR1_BIT_DONE_D2_PT_0
    );
  UAR1_BIT_DONE_D2_107 : X_OR2 
    port map (
      I0 => UAR1_BIT_DONE_D2_PT_0,
      I1 => UAR1_BIT_DONE_D2_PT_0,
      O => UAR1_BIT_DONE_D2
    );
  UAR1_BIT_DONE_XOR : X_XOR2 
    port map (
      I0 => UAR1_BIT_DONE_D1,
      I1 => UAR1_BIT_DONE_D2,
      O => UAR1_BIT_DONE_D
    );
  UAR1_BIT_DONE_FBK_108 : X_BUF 
    port map (
      I => UAR1_BIT_DONE_Q,
      O => UAR1_BIT_DONE_FBK
    );
  UAR1_BC1_CURRENT_STATE_11_Q_109 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_Q,
      O => UAR1_BC1_CURRENT_STATE_11_Q_5
    );
  UAR1_BC1_CURRENT_STATE_11_REG : X_FF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => FSRIO_0,
      RST => PRLD,
      O => UAR1_BC1_CURRENT_STATE_11_Q
    );
  UAR1_BC1_CURRENT_STATE_11_D1_110 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BC1_CURRENT_STATE_11_D1
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_0_111 : X_AND2 
    port map (
      I0 => EXP9_EXP,
      I1 => EXP9_EXP,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_0
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_1_112 : X_AND2 
    port map (
      I0 => EXP10_EXP,
      I1 => EXP10_EXP,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_1
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_2_113 : X_AND7 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_11_D2_PT_2_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_3_FBK,
      I2 => UAR1_BC1_CURRENT_STATE_11_D2_PT_2_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_11_D2_PT_2_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_11_D2_PT_2_4_INV,
      I5 => UAR1_BC1_CURRENT_STATE_11_D2_PT_2_5_INV,
      I6 => UAR1_BC1_CURRENT_STATE_11_D2_PT_2_6_INV,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_2
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_3_114 : X_AND7 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_11_D2_PT_3_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_11_D2_PT_3_1_INV,
      I2 => UAR1_BC1_CURRENT_STATE_11_D2_PT_3_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_11_D2_PT_3_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_2_FBK,
      I5 => UAR1_BC1_CURRENT_STATE_11_D2_PT_3_5_INV,
      I6 => UAR1_BC1_CURRENT_STATE_11_D2_PT_3_6_INV,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_3
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_4_115 : X_AND7 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_11_D2_PT_4_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_11_D2_PT_4_1_INV,
      I2 => UAR1_BC1_CURRENT_STATE_11_D2_PT_4_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_11_D2_PT_4_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_6_FBK,
      I5 => UAR1_BC1_CURRENT_STATE_11_D2_PT_4_5_INV,
      I6 => UAR1_BC1_CURRENT_STATE_11_D2_PT_4_6_INV,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_4
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_5_116 : X_AND7 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_11_D2_PT_5_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_11_D2_PT_5_1_INV,
      I2 => UAR1_BC1_CURRENT_STATE_11_D2_PT_5_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_11_D2_PT_5_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_7_FBK,
      I5 => UAR1_BC1_CURRENT_STATE_11_D2_PT_5_5_INV,
      I6 => UAR1_BC1_CURRENT_STATE_11_D2_PT_5_6_INV,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_5
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_6_117 : X_AND7 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_11_D2_PT_6_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_11_D2_PT_6_1_INV,
      I2 => UAR1_BC1_CURRENT_STATE_11_D2_PT_6_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_11_D2_PT_6_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_8_FBK,
      I5 => UAR1_BC1_CURRENT_STATE_11_D2_PT_6_5_INV,
      I6 => UAR1_BC1_CURRENT_STATE_11_D2_PT_6_6_INV,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_6
    );
  UAR1_BC1_CURRENT_STATE_11_D2_118 : X_OR7 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_11_D2_PT_0,
      I1 => UAR1_BC1_CURRENT_STATE_11_D2_PT_1,
      I2 => UAR1_BC1_CURRENT_STATE_11_D2_PT_2,
      I3 => UAR1_BC1_CURRENT_STATE_11_D2_PT_3,
      I4 => UAR1_BC1_CURRENT_STATE_11_D2_PT_4,
      I5 => UAR1_BC1_CURRENT_STATE_11_D2_PT_5,
      I6 => UAR1_BC1_CURRENT_STATE_11_D2_PT_6,
      O => UAR1_BC1_CURRENT_STATE_11_D2
    );
  UAR1_BC1_CURRENT_STATE_11_XOR : X_XOR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_11_XOR_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_11_D2,
      O => UAR1_BC1_CURRENT_STATE_11_D
    );
  UAR1_BC1_CURRENT_STATE_11_FBK_119 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_Q,
      O => UAR1_BC1_CURRENT_STATE_11_FBK
    );
  EXP9_EXP_PT_0_120 : X_AND6 
    port map (
      I0 => UAR1_DATA_IN,
      I1 => EXP9_EXP_PT_0_1_INV,
      I2 => UAR1_BM1_SAMPLED_BITS(0),
      I3 => UAR1_BM1_SAMPLED_BITS(1),
      I4 => UAR1_BM1_SAMPLED_BITS(2),
      I5 => EXP9_EXP_PT_0_5_INV,
      O => EXP9_EXP_PT_0
    );
  EXP9_EXP_PT_1_121 : X_AND6 
    port map (
      I0 => UAR1_DATA_IN,
      I1 => EXP9_EXP_PT_1_1_INV,
      I2 => EXP9_EXP_PT_1_2_INV,
      I3 => EXP9_EXP_PT_1_3_INV,
      I4 => EXP9_EXP_PT_1_4_INV,
      I5 => EXP9_EXP_PT_1_5_INV,
      O => EXP9_EXP_PT_1
    );
  EXP9_EXP_PT_2_122 : X_AND6 
    port map (
      I0 => EXP9_EXP_PT_2_0_INV,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => EXP9_EXP_PT_2_4_INV,
      I5 => EXP9_EXP_PT_2_5_INV,
      O => EXP9_EXP_PT_2
    );
  EXP9_EXP_PT_3_123 : X_AND7 
    port map (
      I0 => EXP9_EXP_PT_3_0_INV,
      I1 => EXP9_EXP_PT_3_1_INV,
      I2 => EXP9_EXP_PT_3_2_INV,
      I3 => EXP9_EXP_PT_3_3_INV,
      I4 => EXP9_EXP_PT_3_4_INV,
      I5 => UAR1_BC1_CURRENT_STATE_1_FBK,
      I6 => EXP9_EXP_PT_3_6_INV,
      O => EXP9_EXP_PT_3
    );
  EXP9_EXP_PT_4_124 : X_AND16 
    port map (
      I0 => UAR1_DATA_IN,
      I1 => EXP9_EXP_PT_4_1_INV,
      I2 => EXP9_EXP_PT_4_2_INV,
      I3 => EXP9_EXP_PT_4_3_INV,
      I4 => EXP9_EXP_PT_4_4_INV,
      I5 => EXP9_EXP_PT_4_5_INV,
      I6 => EXP9_EXP_PT_4_6_INV,
      I7 => EXP9_EXP_PT_4_7_INV,
      I8 => EXP9_EXP_PT_4_8_INV,
      I9 => EXP9_EXP_PT_4_9_INV,
      I10 => EXP9_EXP_PT_4_10_INV,
      I11 => EXP9_EXP_PT_4_11_INV,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP9_EXP_PT_4
    );
  EXP9_EXP_125 : X_OR5 
    port map (
      I0 => EXP9_EXP_PT_0,
      I1 => EXP9_EXP_PT_1,
      I2 => EXP9_EXP_PT_2,
      I3 => EXP9_EXP_PT_3,
      I4 => EXP9_EXP_PT_4,
      O => EXP9_EXP
    );
  UAR1_DATA_IN_126 : X_BUF 
    port map (
      I => UAR1_DATA_IN_Q,
      O => UAR1_DATA_IN
    );
  UAR1_DATA_IN_R_OR_PRLD_127 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_DATA_IN_R_OR_PRLD
    );
  UAR1_DATA_IN_REG : X_FF 
    port map (
      I => UAR1_DATA_IN_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_DATA_IN_R_OR_PRLD,
      O => UAR1_DATA_IN_Q
    );
  UAR1_DATA_IN_D1_128 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_DATA_IN_D1
    );
  UAR1_DATA_IN_D2_PT_0_129 : X_AND2 
    port map (
      I0 => IR_DETECT_C,
      I1 => IR_DETECT_C,
      O => UAR1_DATA_IN_D2_PT_0
    );
  UAR1_DATA_IN_D2_130 : X_OR2 
    port map (
      I0 => UAR1_DATA_IN_D2_PT_0,
      I1 => UAR1_DATA_IN_D2_PT_0,
      O => UAR1_DATA_IN_D2
    );
  UAR1_DATA_IN_XOR : X_XOR2 
    port map (
      I0 => UAR1_DATA_IN_D1,
      I1 => UAR1_DATA_IN_D2,
      O => UAR1_DATA_IN_D
    );
  UAR1_DATA_IN_FBK_131 : X_BUF 
    port map (
      I => UAR1_DATA_IN_Q,
      O => UAR1_DATA_IN_FBK
    );
  IR_DETECT_C_132 : X_BUF 
    port map (
      I => IR_DETECT,
      O => IR_DETECT_C
    );
  CLK_C_FCLK_133 : X_BUF 
    port map (
      I => CLK,
      O => CLK_C_FCLK
    );
  RESET_C_134 : X_BUF 
    port map (
      I => RESET,
      O => RESET_C
    );
  FSRIO_0_135 : X_BUF 
    port map (
      I => RESET,
      O => FSRIO_0
    );
  UAR1_BM1_SAMPLED_BITS_0_Q_136 : X_BUF 
    port map (
      I => UAR1_BM1_SAMPLED_BITS_0_Q,
      O => UAR1_BM1_SAMPLED_BITS(0)
    );
  UAR1_BM1_SAMPLED_BITS_0_R_OR_PRLD_137 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BM1_SAMPLED_BITS_0_R_OR_PRLD
    );
  UAR1_BM1_SAMPLED_BITS_0_REG : X_FF 
    port map (
      I => UAR1_BM1_SAMPLED_BITS_0_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BM1_SAMPLED_BITS_0_R_OR_PRLD,
      O => UAR1_BM1_SAMPLED_BITS_0_Q
    );
  UAR1_BM1_SAMPLED_BITS_0_D1_138 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BM1_SAMPLED_BITS_0_D1
    );
  UAR1_BM1_SAMPLED_BITS_0_D2_PT_0_139 : X_AND2 
    port map (
      I0 => UAR1_DATA_IN_FBK,
      I1 => UAR1_BM1_CURRENT_STATE_3_FBK,
      O => UAR1_BM1_SAMPLED_BITS_0_D2_PT_0
    );
  UAR1_BM1_SAMPLED_BITS_0_D2_PT_1_140 : X_AND2 
    port map (
      I0 => UAR1_BM1_SAMPLED_BITS_0_D2_PT_1_0_INV,
      I1 => UAR1_BM1_SAMPLED_BITS_0_FBK,
      O => UAR1_BM1_SAMPLED_BITS_0_D2_PT_1
    );
  UAR1_BM1_SAMPLED_BITS_0_D2_141 : X_OR2 
    port map (
      I0 => UAR1_BM1_SAMPLED_BITS_0_D2_PT_0,
      I1 => UAR1_BM1_SAMPLED_BITS_0_D2_PT_1,
      O => UAR1_BM1_SAMPLED_BITS_0_D2
    );
  UAR1_BM1_SAMPLED_BITS_0_XOR : X_XOR2 
    port map (
      I0 => UAR1_BM1_SAMPLED_BITS_0_D1,
      I1 => UAR1_BM1_SAMPLED_BITS_0_D2,
      O => UAR1_BM1_SAMPLED_BITS_0_D
    );
  UAR1_BM1_SAMPLED_BITS_0_FBK_142 : X_BUF 
    port map (
      I => UAR1_BM1_SAMPLED_BITS_0_Q,
      O => UAR1_BM1_SAMPLED_BITS_0_FBK
    );
  UAR1_BM1_CURRENT_STATE_3_FBK_143 : X_BUF 
    port map (
      I => UAR1_BM1_CURRENT_STATE_3_Q,
      O => UAR1_BM1_CURRENT_STATE_3_FBK
    );
  UAR1_BM1_CURRENT_STATE_3_R_OR_PRLD_144 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BM1_CURRENT_STATE_3_R_OR_PRLD
    );
  UAR1_BM1_CURRENT_STATE_3_REG : X_FF 
    port map (
      I => UAR1_BM1_CURRENT_STATE_3_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BM1_CURRENT_STATE_3_R_OR_PRLD,
      O => UAR1_BM1_CURRENT_STATE_3_Q
    );
  UAR1_BM1_CURRENT_STATE_3_D1_145 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BM1_CURRENT_STATE_3_D1
    );
  UAR1_BM1_CURRENT_STATE_3_D2_PT_0_146 : X_AND3 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_3_D2_PT_0_0_INV,
      I1 => UAR1_BM1_CURRENT_STATE_3_D2_PT_0_1_INV,
      I2 => UAR1_BIT_DONE_FBK,
      O => UAR1_BM1_CURRENT_STATE_3_D2_PT_0
    );
  UAR1_BM1_CURRENT_STATE_3_D2_PT_1_147 : X_AND3 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_3_D2_PT_1_0_INV,
      I1 => UAR1_DATA_IN_FBK,
      I2 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_FBK,
      O => UAR1_BM1_CURRENT_STATE_3_D2_PT_1
    );
  UAR1_BM1_CURRENT_STATE_3_D2_148 : X_OR2 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_3_D2_PT_0,
      I1 => UAR1_BM1_CURRENT_STATE_3_D2_PT_1,
      O => UAR1_BM1_CURRENT_STATE_3_D2
    );
  UAR1_BM1_CURRENT_STATE_3_XOR : X_XOR2 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_3_D1,
      I1 => UAR1_BM1_CURRENT_STATE_3_D2,
      O => UAR1_BM1_CURRENT_STATE_3_D
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_FBK_149 : X_BUF 
    port map (
      I => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_Q,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_FBK
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_REG : X_FF 
    port map (
      I => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => FSRIO_0,
      RST => PRLD,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_Q
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D1_150 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D1
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_0_151 : X_AND3 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_0_0_INV,
      I1 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_0_1_INV,
      I2 => UAR1_DATA_IN_FBK,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_0
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_152 : X_AND3 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_0_INV,
      I1 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_1_INV,
      I2 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_2_INV,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_153 : X_AND5 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_0_INV,
      I1 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_1_INV,
      I2 => UAR1_DATA_IN_FBK,
      I3 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_3_INV,
      I4 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_4_INV,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_154 : X_OR3 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_0,
      I1 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1,
      I2 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_XOR : X_XOR2 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_XOR_0_INV,
      I1 => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D
    );
  UAR1_BM1_CURRENT_STATE_1_FBK_155 : X_BUF 
    port map (
      I => UAR1_BM1_CURRENT_STATE_1_Q,
      O => UAR1_BM1_CURRENT_STATE_1_FBK
    );
  UAR1_BM1_CURRENT_STATE_1_R_OR_PRLD_156 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BM1_CURRENT_STATE_1_R_OR_PRLD
    );
  UAR1_BM1_CURRENT_STATE_1_REG : X_FF 
    port map (
      I => UAR1_BM1_CURRENT_STATE_1_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BM1_CURRENT_STATE_1_R_OR_PRLD,
      O => UAR1_BM1_CURRENT_STATE_1_Q
    );
  UAR1_BM1_CURRENT_STATE_1_D1_157 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BM1_CURRENT_STATE_1_D1
    );
  UAR1_BM1_CURRENT_STATE_1_D2_PT_0_158 : X_AND3 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_1_D2_PT_0_0_INV,
      I1 => UAR1_BM1_CURRENT_STATE_1_D2_PT_0_1_INV,
      I2 => UAR1_BM1_CURRENT_STATE_2_FBK,
      O => UAR1_BM1_CURRENT_STATE_1_D2_PT_0
    );
  UAR1_BM1_CURRENT_STATE_1_D2_159 : X_OR2 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_1_D2_PT_0,
      I1 => UAR1_BM1_CURRENT_STATE_1_D2_PT_0,
      O => UAR1_BM1_CURRENT_STATE_1_D2
    );
  UAR1_BM1_CURRENT_STATE_1_XOR : X_XOR2 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_1_D1,
      I1 => UAR1_BM1_CURRENT_STATE_1_D2,
      O => UAR1_BM1_CURRENT_STATE_1_D
    );
  UAR1_BM1_CURRENT_STATE_2_FBK_160 : X_BUF 
    port map (
      I => UAR1_BM1_CURRENT_STATE_2_Q,
      O => UAR1_BM1_CURRENT_STATE_2_FBK
    );
  UAR1_BM1_CURRENT_STATE_2_R_OR_PRLD_161 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BM1_CURRENT_STATE_2_R_OR_PRLD
    );
  UAR1_BM1_CURRENT_STATE_2_REG : X_FF 
    port map (
      I => UAR1_BM1_CURRENT_STATE_2_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BM1_CURRENT_STATE_2_R_OR_PRLD,
      O => UAR1_BM1_CURRENT_STATE_2_Q
    );
  UAR1_BM1_CURRENT_STATE_2_D1_162 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BM1_CURRENT_STATE_2_D1
    );
  UAR1_BM1_CURRENT_STATE_2_D2_PT_0_163 : X_AND3 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_2_D2_PT_0_0_INV,
      I1 => UAR1_BM1_CURRENT_STATE_2_D2_PT_0_1_INV,
      I2 => UAR1_BM1_CURRENT_STATE_3_FBK,
      O => UAR1_BM1_CURRENT_STATE_2_D2_PT_0
    );
  UAR1_BM1_CURRENT_STATE_2_D2_164 : X_OR2 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_2_D2_PT_0,
      I1 => UAR1_BM1_CURRENT_STATE_2_D2_PT_0,
      O => UAR1_BM1_CURRENT_STATE_2_D2
    );
  UAR1_BM1_CURRENT_STATE_2_XOR : X_XOR2 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_2_D1,
      I1 => UAR1_BM1_CURRENT_STATE_2_D2,
      O => UAR1_BM1_CURRENT_STATE_2_D
    );
  UAR1_BM1_SAMPLED_BITS_1_Q_165 : X_BUF 
    port map (
      I => UAR1_BM1_SAMPLED_BITS_1_Q,
      O => UAR1_BM1_SAMPLED_BITS(1)
    );
  UAR1_BM1_SAMPLED_BITS_1_R_OR_PRLD_166 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BM1_SAMPLED_BITS_1_R_OR_PRLD
    );
  UAR1_BM1_SAMPLED_BITS_1_REG : X_FF 
    port map (
      I => UAR1_BM1_SAMPLED_BITS_1_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BM1_SAMPLED_BITS_1_R_OR_PRLD,
      O => UAR1_BM1_SAMPLED_BITS_1_Q
    );
  UAR1_BM1_SAMPLED_BITS_1_D1_167 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BM1_SAMPLED_BITS_1_D1
    );
  UAR1_BM1_SAMPLED_BITS_1_D2_PT_0_168 : X_AND2 
    port map (
      I0 => UAR1_DATA_IN_FBK,
      I1 => UAR1_BM1_CURRENT_STATE_2_FBK,
      O => UAR1_BM1_SAMPLED_BITS_1_D2_PT_0
    );
  UAR1_BM1_SAMPLED_BITS_1_D2_PT_1_169 : X_AND2 
    port map (
      I0 => UAR1_BM1_SAMPLED_BITS_1_D2_PT_1_0_INV,
      I1 => UAR1_BM1_SAMPLED_BITS_1_FBK,
      O => UAR1_BM1_SAMPLED_BITS_1_D2_PT_1
    );
  UAR1_BM1_SAMPLED_BITS_1_D2_170 : X_OR2 
    port map (
      I0 => UAR1_BM1_SAMPLED_BITS_1_D2_PT_0,
      I1 => UAR1_BM1_SAMPLED_BITS_1_D2_PT_1,
      O => UAR1_BM1_SAMPLED_BITS_1_D2
    );
  UAR1_BM1_SAMPLED_BITS_1_XOR : X_XOR2 
    port map (
      I0 => UAR1_BM1_SAMPLED_BITS_1_D1,
      I1 => UAR1_BM1_SAMPLED_BITS_1_D2,
      O => UAR1_BM1_SAMPLED_BITS_1_D
    );
  UAR1_BM1_SAMPLED_BITS_1_FBK_171 : X_BUF 
    port map (
      I => UAR1_BM1_SAMPLED_BITS_1_Q,
      O => UAR1_BM1_SAMPLED_BITS_1_FBK
    );
  UAR1_BM1_SAMPLED_BITS_2_Q_172 : X_BUF 
    port map (
      I => UAR1_BM1_SAMPLED_BITS_2_Q,
      O => UAR1_BM1_SAMPLED_BITS(2)
    );
  UAR1_BM1_SAMPLED_BITS_2_R_OR_PRLD_173 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BM1_SAMPLED_BITS_2_R_OR_PRLD
    );
  UAR1_BM1_SAMPLED_BITS_2_REG : X_FF 
    port map (
      I => UAR1_BM1_SAMPLED_BITS_2_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BM1_SAMPLED_BITS_2_R_OR_PRLD,
      O => UAR1_BM1_SAMPLED_BITS_2_Q
    );
  UAR1_BM1_SAMPLED_BITS_2_D1_174 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BM1_SAMPLED_BITS_2_D1
    );
  UAR1_BM1_SAMPLED_BITS_2_D2_PT_0_175 : X_AND2 
    port map (
      I0 => UAR1_BM1_CURRENT_STATE_1_FBK,
      I1 => UAR1_DATA_IN_FBK,
      O => UAR1_BM1_SAMPLED_BITS_2_D2_PT_0
    );
  UAR1_BM1_SAMPLED_BITS_2_D2_PT_1_176 : X_AND2 
    port map (
      I0 => UAR1_BM1_SAMPLED_BITS_2_D2_PT_1_0_INV,
      I1 => UAR1_BM1_SAMPLED_BITS_2_FBK,
      O => UAR1_BM1_SAMPLED_BITS_2_D2_PT_1
    );
  UAR1_BM1_SAMPLED_BITS_2_D2_177 : X_OR2 
    port map (
      I0 => UAR1_BM1_SAMPLED_BITS_2_D2_PT_0,
      I1 => UAR1_BM1_SAMPLED_BITS_2_D2_PT_1,
      O => UAR1_BM1_SAMPLED_BITS_2_D2
    );
  UAR1_BM1_SAMPLED_BITS_2_XOR : X_XOR2 
    port map (
      I0 => UAR1_BM1_SAMPLED_BITS_2_D1,
      I1 => UAR1_BM1_SAMPLED_BITS_2_D2,
      O => UAR1_BM1_SAMPLED_BITS_2_D
    );
  UAR1_BM1_SAMPLED_BITS_2_FBK_178 : X_BUF 
    port map (
      I => UAR1_BM1_SAMPLED_BITS_2_Q,
      O => UAR1_BM1_SAMPLED_BITS_2_FBK
    );
  UAR1_BC1_CURRENT_STATE_1_Q_179 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_1_Q,
      O => UAR1_BC1_CURRENT_STATE_1_Q_4
    );
  UAR1_BC1_CURRENT_STATE_1_R_OR_PRLD_180 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BC1_CURRENT_STATE_1_R_OR_PRLD
    );
  UAR1_BC1_CURRENT_STATE_1_REG : X_FF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_1_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BC1_CURRENT_STATE_1_R_OR_PRLD,
      O => UAR1_BC1_CURRENT_STATE_1_Q
    );
  UAR1_BC1_CURRENT_STATE_1_D1_181 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BC1_CURRENT_STATE_1_D1
    );
  UAR1_BC1_CURRENT_STATE_1_D2_PT_0_182 : X_AND2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_1_D2_PT_0_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_1_FBK,
      O => UAR1_BC1_CURRENT_STATE_1_D2_PT_0
    );
  UAR1_BC1_CURRENT_STATE_1_D2_PT_1_183 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_2_FBK,
      O => UAR1_BC1_CURRENT_STATE_1_D2_PT_1
    );
  UAR1_BC1_CURRENT_STATE_1_D2_PT_2_184 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BC1_CURRENT_STATE_1_D2_PT_2_1_INV,
      I2 => UAR1_BC1_CURRENT_STATE_1_D2_PT_2_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_1_D2_PT_2_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_2_FBK,
      O => UAR1_BC1_CURRENT_STATE_1_D2_PT_2
    );
  UAR1_BC1_CURRENT_STATE_1_D2_185 : X_OR3 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_1_D2_PT_0,
      I1 => UAR1_BC1_CURRENT_STATE_1_D2_PT_1,
      I2 => UAR1_BC1_CURRENT_STATE_1_D2_PT_2,
      O => UAR1_BC1_CURRENT_STATE_1_D2
    );
  UAR1_BC1_CURRENT_STATE_1_XOR : X_XOR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_1_D1,
      I1 => UAR1_BC1_CURRENT_STATE_1_D2,
      O => UAR1_BC1_CURRENT_STATE_1_D
    );
  UAR1_BC1_CURRENT_STATE_1_FBK_186 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_1_Q,
      O => UAR1_BC1_CURRENT_STATE_1_FBK
    );
  UAR1_BC1_CURRENT_STATE_2_Q_187 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_2_Q,
      O => UAR1_BC1_CURRENT_STATE_2_Q_7
    );
  UAR1_BC1_CURRENT_STATE_2_R_OR_PRLD_188 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BC1_CURRENT_STATE_2_R_OR_PRLD
    );
  UAR1_BC1_CURRENT_STATE_2_REG : X_FF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_2_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BC1_CURRENT_STATE_2_R_OR_PRLD,
      O => UAR1_BC1_CURRENT_STATE_2_Q
    );
  UAR1_BC1_CURRENT_STATE_2_D1_189 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BC1_CURRENT_STATE_2_D1
    );
  UAR1_BC1_CURRENT_STATE_2_D2_PT_0_190 : X_AND2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_2_D2_PT_0_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_2_FBK,
      O => UAR1_BC1_CURRENT_STATE_2_D2_PT_0
    );
  UAR1_BC1_CURRENT_STATE_2_D2_PT_1_191 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BC1_CURRENT_STATE_3_FBK,
      I2 => UAR1_BM1_SAMPLED_BITS(0),
      I3 => UAR1_BM1_SAMPLED_BITS(1),
      I4 => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_2_D2_PT_1
    );
  UAR1_BC1_CURRENT_STATE_2_D2_PT_2_192 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BC1_CURRENT_STATE_3_FBK,
      I2 => UAR1_BC1_CURRENT_STATE_2_D2_PT_2_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_2_D2_PT_2_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_2_D2_PT_2_4_INV,
      O => UAR1_BC1_CURRENT_STATE_2_D2_PT_2
    );
  UAR1_BC1_CURRENT_STATE_2_D2_193 : X_OR3 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_2_D2_PT_0,
      I1 => UAR1_BC1_CURRENT_STATE_2_D2_PT_1,
      I2 => UAR1_BC1_CURRENT_STATE_2_D2_PT_2,
      O => UAR1_BC1_CURRENT_STATE_2_D2
    );
  UAR1_BC1_CURRENT_STATE_2_XOR : X_XOR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_2_D1,
      I1 => UAR1_BC1_CURRENT_STATE_2_D2,
      O => UAR1_BC1_CURRENT_STATE_2_D
    );
  UAR1_BC1_CURRENT_STATE_2_FBK_194 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_2_Q,
      O => UAR1_BC1_CURRENT_STATE_2_FBK
    );
  UAR1_BC1_CURRENT_STATE_3_Q_195 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_3_Q,
      O => UAR1_BC1_CURRENT_STATE_3_Q_8
    );
  UAR1_BC1_CURRENT_STATE_3_R_OR_PRLD_196 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BC1_CURRENT_STATE_3_R_OR_PRLD
    );
  UAR1_BC1_CURRENT_STATE_3_REG : X_FF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_3_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BC1_CURRENT_STATE_3_R_OR_PRLD,
      O => UAR1_BC1_CURRENT_STATE_3_Q
    );
  UAR1_BC1_CURRENT_STATE_3_D1_197 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BC1_CURRENT_STATE_3_D1
    );
  UAR1_BC1_CURRENT_STATE_3_D2_PT_0_198 : X_AND2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_3_D2_PT_0_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_3_FBK,
      O => UAR1_BC1_CURRENT_STATE_3_D2_PT_0
    );
  UAR1_BC1_CURRENT_STATE_3_D2_PT_1_199 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_4_FBK,
      O => UAR1_BC1_CURRENT_STATE_3_D2_PT_1
    );
  UAR1_BC1_CURRENT_STATE_3_D2_PT_2_200 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BC1_CURRENT_STATE_3_D2_PT_2_1_INV,
      I2 => UAR1_BC1_CURRENT_STATE_3_D2_PT_2_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_3_D2_PT_2_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_4_FBK,
      O => UAR1_BC1_CURRENT_STATE_3_D2_PT_2
    );
  UAR1_BC1_CURRENT_STATE_3_D2_201 : X_OR3 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_3_D2_PT_0,
      I1 => UAR1_BC1_CURRENT_STATE_3_D2_PT_1,
      I2 => UAR1_BC1_CURRENT_STATE_3_D2_PT_2,
      O => UAR1_BC1_CURRENT_STATE_3_D2
    );
  UAR1_BC1_CURRENT_STATE_3_XOR : X_XOR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_3_D1,
      I1 => UAR1_BC1_CURRENT_STATE_3_D2,
      O => UAR1_BC1_CURRENT_STATE_3_D
    );
  UAR1_BC1_CURRENT_STATE_3_FBK_202 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_3_Q,
      O => UAR1_BC1_CURRENT_STATE_3_FBK
    );
  UAR1_BC1_CURRENT_STATE_4_FBK_203 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_4_Q,
      O => UAR1_BC1_CURRENT_STATE_4_FBK
    );
  UAR1_BC1_CURRENT_STATE_4_R_OR_PRLD_204 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BC1_CURRENT_STATE_4_R_OR_PRLD
    );
  UAR1_BC1_CURRENT_STATE_4_REG : X_FF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_4_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BC1_CURRENT_STATE_4_R_OR_PRLD,
      O => UAR1_BC1_CURRENT_STATE_4_Q
    );
  UAR1_BC1_CURRENT_STATE_4_D1_205 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BC1_CURRENT_STATE_4_D1
    );
  UAR1_BC1_CURRENT_STATE_4_D2_PT_0_206 : X_AND2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_4_D2_PT_0_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_4_FBK,
      O => UAR1_BC1_CURRENT_STATE_4_D2_PT_0
    );
  UAR1_BC1_CURRENT_STATE_4_D2_PT_1_207 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_5_FBK,
      O => UAR1_BC1_CURRENT_STATE_4_D2_PT_1
    );
  UAR1_BC1_CURRENT_STATE_4_D2_PT_2_208 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BC1_CURRENT_STATE_4_D2_PT_2_1_INV,
      I2 => UAR1_BC1_CURRENT_STATE_4_D2_PT_2_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_4_D2_PT_2_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_5_FBK,
      O => UAR1_BC1_CURRENT_STATE_4_D2_PT_2
    );
  UAR1_BC1_CURRENT_STATE_4_D2_209 : X_OR3 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_4_D2_PT_0,
      I1 => UAR1_BC1_CURRENT_STATE_4_D2_PT_1,
      I2 => UAR1_BC1_CURRENT_STATE_4_D2_PT_2,
      O => UAR1_BC1_CURRENT_STATE_4_D2
    );
  UAR1_BC1_CURRENT_STATE_4_XOR : X_XOR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_4_D1,
      I1 => UAR1_BC1_CURRENT_STATE_4_D2,
      O => UAR1_BC1_CURRENT_STATE_4_D
    );
  UAR1_BC1_CURRENT_STATE_5_FBK_210 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_5_Q,
      O => UAR1_BC1_CURRENT_STATE_5_FBK
    );
  UAR1_BC1_CURRENT_STATE_5_R_OR_PRLD_211 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BC1_CURRENT_STATE_5_R_OR_PRLD
    );
  UAR1_BC1_CURRENT_STATE_5_REG : X_FF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_5_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BC1_CURRENT_STATE_5_R_OR_PRLD,
      O => UAR1_BC1_CURRENT_STATE_5_Q
    );
  UAR1_BC1_CURRENT_STATE_5_D1_212 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BC1_CURRENT_STATE_5_D1
    );
  UAR1_BC1_CURRENT_STATE_5_D2_PT_0_213 : X_AND2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_5_D2_PT_0_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_5_FBK,
      O => UAR1_BC1_CURRENT_STATE_5_D2_PT_0
    );
  UAR1_BC1_CURRENT_STATE_5_D2_PT_1_214 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_6_FBK,
      O => UAR1_BC1_CURRENT_STATE_5_D2_PT_1
    );
  UAR1_BC1_CURRENT_STATE_5_D2_PT_2_215 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BC1_CURRENT_STATE_5_D2_PT_2_1_INV,
      I2 => UAR1_BC1_CURRENT_STATE_5_D2_PT_2_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_5_D2_PT_2_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_6_FBK,
      O => UAR1_BC1_CURRENT_STATE_5_D2_PT_2
    );
  UAR1_BC1_CURRENT_STATE_5_D2_216 : X_OR3 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_5_D2_PT_0,
      I1 => UAR1_BC1_CURRENT_STATE_5_D2_PT_1,
      I2 => UAR1_BC1_CURRENT_STATE_5_D2_PT_2,
      O => UAR1_BC1_CURRENT_STATE_5_D2
    );
  UAR1_BC1_CURRENT_STATE_5_XOR : X_XOR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_5_D1,
      I1 => UAR1_BC1_CURRENT_STATE_5_D2,
      O => UAR1_BC1_CURRENT_STATE_5_D
    );
  UAR1_BC1_CURRENT_STATE_6_FBK_217 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_6_Q,
      O => UAR1_BC1_CURRENT_STATE_6_FBK
    );
  UAR1_BC1_CURRENT_STATE_6_R_OR_PRLD_218 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BC1_CURRENT_STATE_6_R_OR_PRLD
    );
  UAR1_BC1_CURRENT_STATE_6_REG : X_FF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_6_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BC1_CURRENT_STATE_6_R_OR_PRLD,
      O => UAR1_BC1_CURRENT_STATE_6_Q
    );
  UAR1_BC1_CURRENT_STATE_6_D1_219 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BC1_CURRENT_STATE_6_D1
    );
  UAR1_BC1_CURRENT_STATE_6_D2_PT_0_220 : X_AND2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_6_D2_PT_0_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_6_FBK,
      O => UAR1_BC1_CURRENT_STATE_6_D2_PT_0
    );
  UAR1_BC1_CURRENT_STATE_6_D2_PT_1_221 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_7_FBK,
      O => UAR1_BC1_CURRENT_STATE_6_D2_PT_1
    );
  UAR1_BC1_CURRENT_STATE_6_D2_PT_2_222 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BC1_CURRENT_STATE_6_D2_PT_2_1_INV,
      I2 => UAR1_BC1_CURRENT_STATE_6_D2_PT_2_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_6_D2_PT_2_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_7_FBK,
      O => UAR1_BC1_CURRENT_STATE_6_D2_PT_2
    );
  UAR1_BC1_CURRENT_STATE_6_D2_223 : X_OR3 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_6_D2_PT_0,
      I1 => UAR1_BC1_CURRENT_STATE_6_D2_PT_1,
      I2 => UAR1_BC1_CURRENT_STATE_6_D2_PT_2,
      O => UAR1_BC1_CURRENT_STATE_6_D2
    );
  UAR1_BC1_CURRENT_STATE_6_XOR : X_XOR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_6_D1,
      I1 => UAR1_BC1_CURRENT_STATE_6_D2,
      O => UAR1_BC1_CURRENT_STATE_6_D
    );
  UAR1_BC1_CURRENT_STATE_7_FBK_224 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_7_Q,
      O => UAR1_BC1_CURRENT_STATE_7_FBK
    );
  UAR1_BC1_CURRENT_STATE_7_R_OR_PRLD_225 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BC1_CURRENT_STATE_7_R_OR_PRLD
    );
  UAR1_BC1_CURRENT_STATE_7_REG : X_FF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_7_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BC1_CURRENT_STATE_7_R_OR_PRLD,
      O => UAR1_BC1_CURRENT_STATE_7_Q
    );
  UAR1_BC1_CURRENT_STATE_7_D1_226 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BC1_CURRENT_STATE_7_D1
    );
  UAR1_BC1_CURRENT_STATE_7_D2_PT_0_227 : X_AND2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_7_D2_PT_0_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_7_FBK,
      O => UAR1_BC1_CURRENT_STATE_7_D2_PT_0
    );
  UAR1_BC1_CURRENT_STATE_7_D2_PT_1_228 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_8_FBK,
      O => UAR1_BC1_CURRENT_STATE_7_D2_PT_1
    );
  UAR1_BC1_CURRENT_STATE_7_D2_PT_2_229 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BC1_CURRENT_STATE_7_D2_PT_2_1_INV,
      I2 => UAR1_BC1_CURRENT_STATE_7_D2_PT_2_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_7_D2_PT_2_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_8_FBK,
      O => UAR1_BC1_CURRENT_STATE_7_D2_PT_2
    );
  UAR1_BC1_CURRENT_STATE_7_D2_230 : X_OR3 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_7_D2_PT_0,
      I1 => UAR1_BC1_CURRENT_STATE_7_D2_PT_1,
      I2 => UAR1_BC1_CURRENT_STATE_7_D2_PT_2,
      O => UAR1_BC1_CURRENT_STATE_7_D2
    );
  UAR1_BC1_CURRENT_STATE_7_XOR : X_XOR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_7_D1,
      I1 => UAR1_BC1_CURRENT_STATE_7_D2,
      O => UAR1_BC1_CURRENT_STATE_7_D
    );
  UAR1_BC1_CURRENT_STATE_8_FBK_231 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_8_Q,
      O => UAR1_BC1_CURRENT_STATE_8_FBK
    );
  UAR1_BC1_CURRENT_STATE_8_R_OR_PRLD_232 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BC1_CURRENT_STATE_8_R_OR_PRLD
    );
  UAR1_BC1_CURRENT_STATE_8_REG : X_FF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_8_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BC1_CURRENT_STATE_8_R_OR_PRLD,
      O => UAR1_BC1_CURRENT_STATE_8_Q
    );
  UAR1_BC1_CURRENT_STATE_8_D1_233 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BC1_CURRENT_STATE_8_D1
    );
  UAR1_BC1_CURRENT_STATE_8_D2_PT_0_234 : X_AND2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_8_D2_PT_0_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_8_FBK,
      O => UAR1_BC1_CURRENT_STATE_8_D2_PT_0
    );
  UAR1_BC1_CURRENT_STATE_8_D2_PT_1_235 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_9_FBK,
      O => UAR1_BC1_CURRENT_STATE_8_D2_PT_1
    );
  UAR1_BC1_CURRENT_STATE_8_D2_PT_2_236 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BC1_CURRENT_STATE_8_D2_PT_2_1_INV,
      I2 => UAR1_BC1_CURRENT_STATE_8_D2_PT_2_2_INV,
      I3 => UAR1_BC1_CURRENT_STATE_8_D2_PT_2_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_9_FBK,
      O => UAR1_BC1_CURRENT_STATE_8_D2_PT_2
    );
  UAR1_BC1_CURRENT_STATE_8_D2_237 : X_OR3 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_8_D2_PT_0,
      I1 => UAR1_BC1_CURRENT_STATE_8_D2_PT_1,
      I2 => UAR1_BC1_CURRENT_STATE_8_D2_PT_2,
      O => UAR1_BC1_CURRENT_STATE_8_D2
    );
  UAR1_BC1_CURRENT_STATE_8_XOR : X_XOR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_8_D1,
      I1 => UAR1_BC1_CURRENT_STATE_8_D2,
      O => UAR1_BC1_CURRENT_STATE_8_D
    );
  UAR1_BC1_CURRENT_STATE_9_FBK_238 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_9_Q,
      O => UAR1_BC1_CURRENT_STATE_9_FBK
    );
  UAR1_BC1_CURRENT_STATE_9_R_OR_PRLD_239 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BC1_CURRENT_STATE_9_R_OR_PRLD
    );
  UAR1_BC1_CURRENT_STATE_9_REG : X_FF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_9_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BC1_CURRENT_STATE_9_R_OR_PRLD,
      O => UAR1_BC1_CURRENT_STATE_9_Q
    );
  UAR1_BC1_CURRENT_STATE_9_D1_240 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BC1_CURRENT_STATE_9_D1
    );
  UAR1_BC1_CURRENT_STATE_9_D2_PT_0_241 : X_AND2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_9_D2_PT_0_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_9_FBK,
      O => UAR1_BC1_CURRENT_STATE_9_D2_PT_0
    );
  UAR1_BC1_CURRENT_STATE_9_D2_PT_1_242 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_10_Q_6,
      O => UAR1_BC1_CURRENT_STATE_9_D2_PT_1
    );
  UAR1_BC1_CURRENT_STATE_9_D2_243 : X_OR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_9_D2_PT_0,
      I1 => UAR1_BC1_CURRENT_STATE_9_D2_PT_1,
      O => UAR1_BC1_CURRENT_STATE_9_D2
    );
  UAR1_BC1_CURRENT_STATE_9_XOR : X_XOR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_9_D1,
      I1 => UAR1_BC1_CURRENT_STATE_9_D2,
      O => UAR1_BC1_CURRENT_STATE_9_D
    );
  UAR1_BC1_CURRENT_STATE_10_Q_244 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q,
      O => UAR1_BC1_CURRENT_STATE_10_Q_6
    );
  UAR1_BC1_CURRENT_STATE_10_R_OR_PRLD_245 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BC1_CURRENT_STATE_10_R_OR_PRLD
    );
  UAR1_BC1_CURRENT_STATE_10_REG : X_FF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BC1_CURRENT_STATE_10_R_OR_PRLD,
      O => UAR1_BC1_CURRENT_STATE_10_Q
    );
  UAR1_BC1_CURRENT_STATE_10_D1_246 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BC1_CURRENT_STATE_10_D1
    );
  UAR1_BC1_CURRENT_STATE_10_D2_PT_0_247 : X_AND2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_11_Q_5,
      I1 => UAR1_DATA_IN_FBK,
      O => UAR1_BC1_CURRENT_STATE_10_D2_PT_0
    );
  UAR1_BC1_CURRENT_STATE_10_D2_PT_1_248 : X_AND2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_10_D2_PT_1_0_INV,
      I1 => UAR1_BC1_CURRENT_STATE_10_FBK,
      O => UAR1_BC1_CURRENT_STATE_10_D2_PT_1
    );
  UAR1_BC1_CURRENT_STATE_10_D2_249 : X_OR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_10_D2_PT_0,
      I1 => UAR1_BC1_CURRENT_STATE_10_D2_PT_1,
      O => UAR1_BC1_CURRENT_STATE_10_D2
    );
  UAR1_BC1_CURRENT_STATE_10_XOR : X_XOR2 
    port map (
      I0 => UAR1_BC1_CURRENT_STATE_10_D1,
      I1 => UAR1_BC1_CURRENT_STATE_10_D2,
      O => UAR1_BC1_CURRENT_STATE_10_D
    );
  UAR1_BC1_CURRENT_STATE_10_FBK_250 : X_BUF 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q,
      O => UAR1_BC1_CURRENT_STATE_10_FBK
    );
  EXP10_EXP_PT_0_251 : X_AND3 
    port map (
      I0 => EXP10_EXP_PT_0_0_INV,
      I1 => UAR1_DATA_IN,
      I2 => EXP10_EXP_PT_0_2_INV,
      O => EXP10_EXP_PT_0
    );
  EXP10_EXP_PT_1_252 : X_AND3 
    port map (
      I0 => EXP10_EXP_PT_1_0_INV,
      I1 => EXP10_EXP_PT_1_1_INV,
      I2 => EXP10_EXP_PT_1_2_INV,
      O => EXP10_EXP_PT_1
    );
  EXP10_EXP_PT_2_253 : X_AND7 
    port map (
      I0 => EXP10_EXP_PT_2_0_INV,
      I1 => EXP10_EXP_PT_2_1_INV,
      I2 => EXP10_EXP_PT_2_2_INV,
      I3 => EXP10_EXP_PT_2_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_4_FBK,
      I5 => EXP10_EXP_PT_2_5_INV,
      I6 => EXP10_EXP_PT_2_6_INV,
      O => EXP10_EXP_PT_2
    );
  EXP10_EXP_PT_3_254 : X_AND7 
    port map (
      I0 => EXP10_EXP_PT_3_0_INV,
      I1 => EXP10_EXP_PT_3_1_INV,
      I2 => EXP10_EXP_PT_3_2_INV,
      I3 => EXP10_EXP_PT_3_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_5_FBK,
      I5 => EXP10_EXP_PT_3_5_INV,
      I6 => EXP10_EXP_PT_3_6_INV,
      O => EXP10_EXP_PT_3
    );
  EXP10_EXP_PT_4_255 : X_AND7 
    port map (
      I0 => EXP10_EXP_PT_4_0_INV,
      I1 => EXP10_EXP_PT_4_1_INV,
      I2 => EXP10_EXP_PT_4_2_INV,
      I3 => EXP10_EXP_PT_4_3_INV,
      I4 => UAR1_BC1_CURRENT_STATE_9_FBK,
      I5 => EXP10_EXP_PT_4_5_INV,
      I6 => EXP10_EXP_PT_4_6_INV,
      O => EXP10_EXP_PT_4
    );
  EXP10_EXP_256 : X_OR5 
    port map (
      I0 => EXP10_EXP_PT_0,
      I1 => EXP10_EXP_PT_1,
      I2 => EXP10_EXP_PT_2,
      I3 => EXP10_EXP_PT_3,
      I4 => EXP10_EXP_PT_4,
      O => EXP10_EXP
    );
  UAR1_BYTE_OUT_7_Q_257 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_7_Q,
      O => UAR1_BYTE_OUT(7)
    );
  UAR1_BYTE_OUT_7_R_OR_PRLD_258 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BYTE_OUT_7_R_OR_PRLD
    );
  UAR1_BYTE_OUT_7_REG : X_FF 
    port map (
      I => UAR1_BYTE_OUT_7_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BYTE_OUT_7_R_OR_PRLD,
      O => UAR1_BYTE_OUT_7_Q
    );
  UAR1_BYTE_OUT_7_D1_259 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BYTE_OUT_7_D1
    );
  UAR1_BYTE_OUT_7_D2_PT_0_260 : X_AND2 
    port map (
      I0 => UAR1_BYTE_OUT_7_D2_PT_0_0_INV,
      I1 => UAR1_BYTE_OUT_7_FBK,
      O => UAR1_BYTE_OUT_7_D2_PT_0
    );
  UAR1_BYTE_OUT_7_D2_PT_1_261 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE_FBK,
      I1 => UAR1_BC1_CURRENT_STATE_2_Q_7,
      I2 => UAR1_BM1_SAMPLED_BITS_0_FBK,
      I3 => UAR1_BM1_SAMPLED_BITS_1_FBK,
      I4 => UAR1_BM1_SAMPLED_BITS_2_FBK,
      O => UAR1_BYTE_OUT_7_D2_PT_1
    );
  UAR1_BYTE_OUT_7_D2_262 : X_OR2 
    port map (
      I0 => UAR1_BYTE_OUT_7_D2_PT_0,
      I1 => UAR1_BYTE_OUT_7_D2_PT_1,
      O => UAR1_BYTE_OUT_7_D2
    );
  UAR1_BYTE_OUT_7_XOR : X_XOR2 
    port map (
      I0 => UAR1_BYTE_OUT_7_D1,
      I1 => UAR1_BYTE_OUT_7_D2,
      O => UAR1_BYTE_OUT_7_D
    );
  UAR1_BYTE_OUT_7_FBK_263 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_7_Q,
      O => UAR1_BYTE_OUT_7_FBK
    );
  RC_ADDRESS_C_1_Q : X_BUF 
    port map (
      I => RC_ADDRESS(1),
      O => RC_ADDRESS_C(1)
    );
  RXD_5_FBK_264 : X_BUF 
    port map (
      I => RXD_5_Q,
      O => RXD_5_FBK
    );
  RXD_5_R_OR_PRLD_265 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => RXD_5_R_OR_PRLD
    );
  RXD_5_REG : X_FF 
    port map (
      I => RXD_5_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => RXD_5_R_OR_PRLD,
      O => RXD_5_Q
    );
  RXD_5_D1_266 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => RXD_5_D1
    );
  RXD_5_D2_PT_0_267 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_5_D2_PT_0_1_INV,
      I2 => RXD_5_FBK,
      I3 => RXD_5_D2_PT_0_3_INV,
      O => RXD_5_D2_PT_0
    );
  RXD_5_D2_PT_1_268 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_5_D2_PT_1_1_INV,
      I2 => RXD_5_D2_PT_1_2_INV,
      I3 => UAR1_BYTE_OUT(5),
      O => RXD_5_D2_PT_1
    );
  RXD_5_D2_269 : X_OR2 
    port map (
      I0 => RXD_5_D2_PT_0,
      I1 => RXD_5_D2_PT_1,
      O => RXD_5_D2
    );
  RXD_5_D_270 : X_XOR2 
    port map (
      I0 => RXD_5_D_TFF,
      I1 => RXD_5_Q,
      O => RXD_5_D
    );
  RXD_5_XOR : X_XOR2 
    port map (
      I0 => RXD_5_D1,
      I1 => RXD_5_D2,
      O => RXD_5_D_TFF
    );
  UAR1_BYTE_OUT_5_Q_271 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_5_Q,
      O => UAR1_BYTE_OUT(5)
    );
  UAR1_BYTE_OUT_5_R_OR_PRLD_272 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BYTE_OUT_5_R_OR_PRLD
    );
  UAR1_BYTE_OUT_5_REG : X_FF 
    port map (
      I => UAR1_BYTE_OUT_5_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BYTE_OUT_5_R_OR_PRLD,
      O => UAR1_BYTE_OUT_5_Q
    );
  UAR1_BYTE_OUT_5_D1_273 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BYTE_OUT_5_D1
    );
  UAR1_BYTE_OUT_5_D2_PT_0_274 : X_AND2 
    port map (
      I0 => UAR1_BYTE_OUT_5_D2_PT_0_0_INV,
      I1 => UAR1_BYTE_OUT_5_FBK,
      O => UAR1_BYTE_OUT_5_D2_PT_0
    );
  UAR1_BYTE_OUT_5_D2_PT_1_275 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_4_FBK,
      O => UAR1_BYTE_OUT_5_D2_PT_1
    );
  UAR1_BYTE_OUT_5_D2_276 : X_OR2 
    port map (
      I0 => UAR1_BYTE_OUT_5_D2_PT_0,
      I1 => UAR1_BYTE_OUT_5_D2_PT_1,
      O => UAR1_BYTE_OUT_5_D2
    );
  UAR1_BYTE_OUT_5_XOR : X_XOR2 
    port map (
      I0 => UAR1_BYTE_OUT_5_D1,
      I1 => UAR1_BYTE_OUT_5_D2,
      O => UAR1_BYTE_OUT_5_D
    );
  UAR1_BYTE_OUT_5_FBK_277 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_5_Q,
      O => UAR1_BYTE_OUT_5_FBK
    );
  RC_ADDRESS_C_2_Q : X_BUF 
    port map (
      I => RC_ADDRESS(2),
      O => RC_ADDRESS_C(2)
    );
  RXD_6_FBK_278 : X_BUF 
    port map (
      I => RXD_6_Q,
      O => RXD_6_FBK
    );
  RXD_6_R_OR_PRLD_279 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => RXD_6_R_OR_PRLD
    );
  RXD_6_REG : X_FF 
    port map (
      I => RXD_6_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => RXD_6_R_OR_PRLD,
      O => RXD_6_Q
    );
  RXD_6_D1_280 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => RXD_6_D1
    );
  RXD_6_D2_PT_0_281 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_6_D2_PT_0_1_INV,
      I2 => RXD_6_FBK,
      I3 => RXD_6_D2_PT_0_3_INV,
      O => RXD_6_D2_PT_0
    );
  RXD_6_D2_PT_1_282 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_6_D2_PT_1_1_INV,
      I2 => RXD_6_D2_PT_1_2_INV,
      I3 => UAR1_BYTE_OUT(6),
      O => RXD_6_D2_PT_1
    );
  RXD_6_D2_283 : X_OR2 
    port map (
      I0 => RXD_6_D2_PT_0,
      I1 => RXD_6_D2_PT_1,
      O => RXD_6_D2
    );
  RXD_6_D_284 : X_XOR2 
    port map (
      I0 => RXD_6_D_TFF,
      I1 => RXD_6_Q,
      O => RXD_6_D
    );
  RXD_6_XOR : X_XOR2 
    port map (
      I0 => RXD_6_D1,
      I1 => RXD_6_D2,
      O => RXD_6_D_TFF
    );
  UAR1_BYTE_OUT_6_Q_285 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_6_Q,
      O => UAR1_BYTE_OUT(6)
    );
  UAR1_BYTE_OUT_6_R_OR_PRLD_286 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BYTE_OUT_6_R_OR_PRLD
    );
  UAR1_BYTE_OUT_6_REG : X_FF 
    port map (
      I => UAR1_BYTE_OUT_6_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BYTE_OUT_6_R_OR_PRLD,
      O => UAR1_BYTE_OUT_6_Q
    );
  UAR1_BYTE_OUT_6_D1_287 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BYTE_OUT_6_D1
    );
  UAR1_BYTE_OUT_6_D2_PT_0_288 : X_AND2 
    port map (
      I0 => UAR1_BYTE_OUT_6_D2_PT_0_0_INV,
      I1 => UAR1_BYTE_OUT_6_FBK,
      O => UAR1_BYTE_OUT_6_D2_PT_0
    );
  UAR1_BYTE_OUT_6_D2_PT_1_289 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE_FBK,
      I1 => UAR1_BC1_CURRENT_STATE_3_Q_8,
      I2 => UAR1_BM1_SAMPLED_BITS_0_FBK,
      I3 => UAR1_BM1_SAMPLED_BITS_1_FBK,
      I4 => UAR1_BM1_SAMPLED_BITS_2_FBK,
      O => UAR1_BYTE_OUT_6_D2_PT_1
    );
  UAR1_BYTE_OUT_6_D2_290 : X_OR2 
    port map (
      I0 => UAR1_BYTE_OUT_6_D2_PT_0,
      I1 => UAR1_BYTE_OUT_6_D2_PT_1,
      O => UAR1_BYTE_OUT_6_D2
    );
  UAR1_BYTE_OUT_6_XOR : X_XOR2 
    port map (
      I0 => UAR1_BYTE_OUT_6_D1,
      I1 => UAR1_BYTE_OUT_6_D2,
      O => UAR1_BYTE_OUT_6_D
    );
  UAR1_BYTE_OUT_6_FBK_291 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_6_Q,
      O => UAR1_BYTE_OUT_6_FBK
    );
  RC_ADDRESS_C_3_Q : X_BUF 
    port map (
      I => RC_ADDRESS(3),
      O => RC_ADDRESS_C(3)
    );
  RXD_2_FBK_292 : X_BUF 
    port map (
      I => RXD_2_Q,
      O => RXD_2_FBK
    );
  RXD_2_R_OR_PRLD_293 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => RXD_2_R_OR_PRLD
    );
  RXD_2_REG : X_FF 
    port map (
      I => RXD_2_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => RXD_2_R_OR_PRLD,
      O => RXD_2_Q
    );
  RXD_2_D1_294 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => RXD_2_D1
    );
  RXD_2_D2_PT_0_295 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_2_D2_PT_0_1_INV,
      I2 => RXD_2_FBK,
      I3 => RXD_2_D2_PT_0_3_INV,
      O => RXD_2_D2_PT_0
    );
  RXD_2_D2_PT_1_296 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_2_D2_PT_1_1_INV,
      I2 => RXD_2_D2_PT_1_2_INV,
      I3 => UAR1_BYTE_OUT(2),
      O => RXD_2_D2_PT_1
    );
  RXD_2_D2_297 : X_OR2 
    port map (
      I0 => RXD_2_D2_PT_0,
      I1 => RXD_2_D2_PT_1,
      O => RXD_2_D2
    );
  RXD_2_D_298 : X_XOR2 
    port map (
      I0 => RXD_2_D_TFF,
      I1 => RXD_2_Q,
      O => RXD_2_D
    );
  RXD_2_XOR : X_XOR2 
    port map (
      I0 => RXD_2_D1,
      I1 => RXD_2_D2,
      O => RXD_2_D_TFF
    );
  UAR1_BYTE_OUT_2_Q_299 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_2_Q,
      O => UAR1_BYTE_OUT(2)
    );
  UAR1_BYTE_OUT_2_R_OR_PRLD_300 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BYTE_OUT_2_R_OR_PRLD
    );
  UAR1_BYTE_OUT_2_REG : X_FF 
    port map (
      I => UAR1_BYTE_OUT_2_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BYTE_OUT_2_R_OR_PRLD,
      O => UAR1_BYTE_OUT_2_Q
    );
  UAR1_BYTE_OUT_2_D1_301 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BYTE_OUT_2_D1
    );
  UAR1_BYTE_OUT_2_D2_PT_0_302 : X_AND2 
    port map (
      I0 => UAR1_BYTE_OUT_2_D2_PT_0_0_INV,
      I1 => UAR1_BYTE_OUT_2_FBK,
      O => UAR1_BYTE_OUT_2_D2_PT_0
    );
  UAR1_BYTE_OUT_2_D2_PT_1_303 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_7_FBK,
      O => UAR1_BYTE_OUT_2_D2_PT_1
    );
  UAR1_BYTE_OUT_2_D2_304 : X_OR2 
    port map (
      I0 => UAR1_BYTE_OUT_2_D2_PT_0,
      I1 => UAR1_BYTE_OUT_2_D2_PT_1,
      O => UAR1_BYTE_OUT_2_D2
    );
  UAR1_BYTE_OUT_2_XOR : X_XOR2 
    port map (
      I0 => UAR1_BYTE_OUT_2_D1,
      I1 => UAR1_BYTE_OUT_2_D2,
      O => UAR1_BYTE_OUT_2_D
    );
  UAR1_BYTE_OUT_2_FBK_305 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_2_Q,
      O => UAR1_BYTE_OUT_2_FBK
    );
  EXP19_EXP_PT_0_306 : X_AND2 
    port map (
      I0 => RC_ADDRESS_C(1),
      I1 => EXP19_EXP_PT_0_1_INV,
      O => EXP19_EXP_PT_0
    );
  EXP19_EXP_PT_1_307 : X_AND2 
    port map (
      I0 => EXP19_EXP_PT_1_0_INV,
      I1 => RXD_5_FBK,
      O => EXP19_EXP_PT_1
    );
  EXP19_EXP_PT_2_308 : X_AND2 
    port map (
      I0 => RC_ADDRESS_C(2),
      I1 => EXP19_EXP_PT_2_1_INV,
      O => EXP19_EXP_PT_2
    );
  EXP19_EXP_PT_3_309 : X_AND2 
    port map (
      I0 => EXP19_EXP_PT_3_0_INV,
      I1 => RXD_6_FBK,
      O => EXP19_EXP_PT_3
    );
  EXP19_EXP_PT_4_310 : X_AND2 
    port map (
      I0 => RC_ADDRESS_C(3),
      I1 => EXP19_EXP_PT_4_1_INV,
      O => EXP19_EXP_PT_4
    );
  EXP19_EXP_311 : X_OR5 
    port map (
      I0 => EXP19_EXP_PT_0,
      I1 => EXP19_EXP_PT_1,
      I2 => EXP19_EXP_PT_2,
      I3 => EXP19_EXP_PT_3,
      I4 => EXP19_EXP_PT_4,
      O => EXP19_EXP
    );
  EXP20_EXP_PT_0_312 : X_AND2 
    port map (
      I0 => RXD_1_EXP,
      I1 => RXD_1_EXP,
      O => EXP20_EXP_PT_0
    );
  EXP20_EXP_PT_1_313 : X_AND2 
    port map (
      I0 => RXD_3_FBK,
      I1 => EXP20_EXP_PT_1_1_INV,
      O => EXP20_EXP_PT_1
    );
  EXP20_EXP_PT_2_314 : X_AND2 
    port map (
      I0 => CM_FADE_DOWN_FBK,
      I1 => RXD_0_FBK,
      O => EXP20_EXP_PT_2
    );
  EXP20_EXP_PT_3_315 : X_AND2 
    port map (
      I0 => EXP20_EXP_PT_3_0_INV,
      I1 => RXD_1_FBK,
      O => EXP20_EXP_PT_3
    );
  EXP20_EXP_PT_4_316 : X_AND2 
    port map (
      I0 => EXP20_EXP_PT_4_0_INV,
      I1 => EXP20_EXP_PT_4_1_INV,
      O => EXP20_EXP_PT_4
    );
  EXP20_EXP_PT_5_317 : X_AND2 
    port map (
      I0 => EXP20_EXP_PT_5_0_INV,
      I1 => RXD_7_FBK,
      O => EXP20_EXP_PT_5
    );
  EXP20_EXP_318 : X_OR6 
    port map (
      I0 => EXP20_EXP_PT_0,
      I1 => EXP20_EXP_PT_1,
      I2 => EXP20_EXP_PT_2,
      I3 => EXP20_EXP_PT_3,
      I4 => EXP20_EXP_PT_4,
      I5 => EXP20_EXP_PT_5,
      O => EXP20_EXP
    );
  RXD_1_EXP_PT_0_319 : X_AND2 
    port map (
      I0 => RXD_3_FBK,
      I1 => RXD_1_FBK,
      O => RXD_1_EXP_PT_0
    );
  RXD_1_EXP_PT_1_320 : X_AND3 
    port map (
      I0 => RXD_1_EXP_PT_1_0_INV,
      I1 => CM_FADE_DOWN_FBK,
      I2 => RXD_1_EXP_PT_1_2_INV,
      O => RXD_1_EXP_PT_1
    );
  RXD_1_EXP_321 : X_OR2 
    port map (
      I0 => RXD_1_EXP_PT_0,
      I1 => RXD_1_EXP_PT_1,
      O => RXD_1_EXP
    );
  RXD_1_FBK_322 : X_BUF 
    port map (
      I => RXD_1_Q,
      O => RXD_1_FBK
    );
  RXD_1_R_OR_PRLD_323 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => RXD_1_R_OR_PRLD
    );
  RXD_1_REG : X_FF 
    port map (
      I => RXD_1_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => RXD_1_R_OR_PRLD,
      O => RXD_1_Q
    );
  RXD_1_D1_324 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => RXD_1_D1
    );
  RXD_1_D2_PT_0_325 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_1_D2_PT_0_1_INV,
      I2 => UAR1_BYTE_OUT(1),
      I3 => RXD_1_D2_PT_0_3_INV,
      O => RXD_1_D2_PT_0
    );
  RXD_1_D2_PT_1_326 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_1_D2_PT_1_1_INV,
      I2 => RXD_1_D2_PT_1_2_INV,
      I3 => RXD_1_FBK,
      O => RXD_1_D2_PT_1
    );
  RXD_1_D2_327 : X_OR2 
    port map (
      I0 => RXD_1_D2_PT_0,
      I1 => RXD_1_D2_PT_1,
      O => RXD_1_D2
    );
  RXD_1_D_328 : X_XOR2 
    port map (
      I0 => RXD_1_D_TFF,
      I1 => RXD_1_Q,
      O => RXD_1_D
    );
  RXD_1_XOR : X_XOR2 
    port map (
      I0 => RXD_1_D1,
      I1 => RXD_1_D2,
      O => RXD_1_D_TFF
    );
  UAR1_BYTE_OUT_1_Q_329 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_1_Q,
      O => UAR1_BYTE_OUT(1)
    );
  UAR1_BYTE_OUT_1_R_OR_PRLD_330 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BYTE_OUT_1_R_OR_PRLD
    );
  UAR1_BYTE_OUT_1_REG : X_FF 
    port map (
      I => UAR1_BYTE_OUT_1_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BYTE_OUT_1_R_OR_PRLD,
      O => UAR1_BYTE_OUT_1_Q
    );
  UAR1_BYTE_OUT_1_D1_331 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BYTE_OUT_1_D1
    );
  UAR1_BYTE_OUT_1_D2_PT_0_332 : X_AND2 
    port map (
      I0 => UAR1_BYTE_OUT_1_D2_PT_0_0_INV,
      I1 => UAR1_BYTE_OUT_1_FBK,
      O => UAR1_BYTE_OUT_1_D2_PT_0
    );
  UAR1_BYTE_OUT_1_D2_PT_1_333 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_8_FBK,
      O => UAR1_BYTE_OUT_1_D2_PT_1
    );
  UAR1_BYTE_OUT_1_D2_334 : X_OR2 
    port map (
      I0 => UAR1_BYTE_OUT_1_D2_PT_0,
      I1 => UAR1_BYTE_OUT_1_D2_PT_1,
      O => UAR1_BYTE_OUT_1_D2
    );
  UAR1_BYTE_OUT_1_XOR : X_XOR2 
    port map (
      I0 => UAR1_BYTE_OUT_1_D1,
      I1 => UAR1_BYTE_OUT_1_D2,
      O => UAR1_BYTE_OUT_1_D
    );
  UAR1_BYTE_OUT_1_FBK_335 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_1_Q,
      O => UAR1_BYTE_OUT_1_FBK
    );
  RXD_3_FBK_336 : X_BUF 
    port map (
      I => RXD_3_Q,
      O => RXD_3_FBK
    );
  RXD_3_R_OR_PRLD_337 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => RXD_3_R_OR_PRLD
    );
  RXD_3_REG : X_FF 
    port map (
      I => RXD_3_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => RXD_3_R_OR_PRLD,
      O => RXD_3_Q
    );
  RXD_3_D1_338 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => RXD_3_D1
    );
  RXD_3_D2_PT_0_339 : X_AND4 
    port map (
      I0 => RXD_3_FBK,
      I1 => UAR1_BYTE_AVAIL,
      I2 => RXD_3_D2_PT_0_2_INV,
      I3 => RXD_3_D2_PT_0_3_INV,
      O => RXD_3_D2_PT_0
    );
  RXD_3_D2_PT_1_340 : X_AND4 
    port map (
      I0 => RXD_3_D2_PT_1_0_INV,
      I1 => UAR1_BYTE_AVAIL,
      I2 => RXD_3_D2_PT_1_2_INV,
      I3 => UAR1_BYTE_OUT(3),
      O => RXD_3_D2_PT_1
    );
  RXD_3_D2_341 : X_OR2 
    port map (
      I0 => RXD_3_D2_PT_0,
      I1 => RXD_3_D2_PT_1,
      O => RXD_3_D2
    );
  RXD_3_D_342 : X_XOR2 
    port map (
      I0 => RXD_3_D_TFF,
      I1 => RXD_3_Q,
      O => RXD_3_D
    );
  RXD_3_XOR : X_XOR2 
    port map (
      I0 => RXD_3_D1,
      I1 => RXD_3_D2,
      O => RXD_3_D_TFF
    );
  UAR1_BYTE_OUT_3_Q_343 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_3_Q,
      O => UAR1_BYTE_OUT(3)
    );
  UAR1_BYTE_OUT_3_R_OR_PRLD_344 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BYTE_OUT_3_R_OR_PRLD
    );
  UAR1_BYTE_OUT_3_REG : X_FF 
    port map (
      I => UAR1_BYTE_OUT_3_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BYTE_OUT_3_R_OR_PRLD,
      O => UAR1_BYTE_OUT_3_Q
    );
  UAR1_BYTE_OUT_3_D1_345 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BYTE_OUT_3_D1
    );
  UAR1_BYTE_OUT_3_D2_PT_0_346 : X_AND2 
    port map (
      I0 => UAR1_BYTE_OUT_3_D2_PT_0_0_INV,
      I1 => UAR1_BYTE_OUT_3_FBK,
      O => UAR1_BYTE_OUT_3_D2_PT_0
    );
  UAR1_BYTE_OUT_3_D2_PT_1_347 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_6_FBK,
      O => UAR1_BYTE_OUT_3_D2_PT_1
    );
  UAR1_BYTE_OUT_3_D2_348 : X_OR2 
    port map (
      I0 => UAR1_BYTE_OUT_3_D2_PT_0,
      I1 => UAR1_BYTE_OUT_3_D2_PT_1,
      O => UAR1_BYTE_OUT_3_D2
    );
  UAR1_BYTE_OUT_3_XOR : X_XOR2 
    port map (
      I0 => UAR1_BYTE_OUT_3_D1,
      I1 => UAR1_BYTE_OUT_3_D2,
      O => UAR1_BYTE_OUT_3_D
    );
  UAR1_BYTE_OUT_3_FBK_349 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_3_Q,
      O => UAR1_BYTE_OUT_3_FBK
    );
  RXD_0_EXP_PT_0_350 : X_AND2 
    port map (
      I0 => RXD_1_FBK,
      I1 => RXD_0_FBK,
      O => RXD_0_EXP_PT_0
    );
  RXD_0_EXP_PT_1_351 : X_AND3 
    port map (
      I0 => RXD_0_EXP_PT_1_0_INV,
      I1 => CM_PANIC_ON_FBK,
      I2 => RXD_0_EXP_PT_1_2_INV,
      O => RXD_0_EXP_PT_1
    );
  RXD_0_EXP_352 : X_OR2 
    port map (
      I0 => RXD_0_EXP_PT_0,
      I1 => RXD_0_EXP_PT_1,
      O => RXD_0_EXP
    );
  RXD_0_FBK_353 : X_BUF 
    port map (
      I => RXD_0_Q,
      O => RXD_0_FBK
    );
  RXD_0_R_OR_PRLD_354 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => RXD_0_R_OR_PRLD
    );
  RXD_0_REG : X_FF 
    port map (
      I => RXD_0_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => RXD_0_R_OR_PRLD,
      O => RXD_0_Q
    );
  RXD_0_D1_355 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => RXD_0_D1
    );
  RXD_0_D2_PT_0_356 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_0_D2_PT_0_1_INV,
      I2 => UAR1_BYTE_OUT(0),
      I3 => RXD_0_D2_PT_0_3_INV,
      O => RXD_0_D2_PT_0
    );
  RXD_0_D2_PT_1_357 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_0_D2_PT_1_1_INV,
      I2 => RXD_0_D2_PT_1_2_INV,
      I3 => RXD_0_FBK,
      O => RXD_0_D2_PT_1
    );
  RXD_0_D2_358 : X_OR2 
    port map (
      I0 => RXD_0_D2_PT_0,
      I1 => RXD_0_D2_PT_1,
      O => RXD_0_D2
    );
  RXD_0_D_359 : X_XOR2 
    port map (
      I0 => RXD_0_D_TFF,
      I1 => RXD_0_Q,
      O => RXD_0_D
    );
  RXD_0_XOR : X_XOR2 
    port map (
      I0 => RXD_0_D1,
      I1 => RXD_0_D2,
      O => RXD_0_D_TFF
    );
  UAR1_BYTE_OUT_0_Q_360 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_0_Q,
      O => UAR1_BYTE_OUT(0)
    );
  UAR1_BYTE_OUT_0_R_OR_PRLD_361 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BYTE_OUT_0_R_OR_PRLD
    );
  UAR1_BYTE_OUT_0_REG : X_FF 
    port map (
      I => UAR1_BYTE_OUT_0_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BYTE_OUT_0_R_OR_PRLD,
      O => UAR1_BYTE_OUT_0_Q
    );
  UAR1_BYTE_OUT_0_D1_362 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BYTE_OUT_0_D1
    );
  UAR1_BYTE_OUT_0_D2_PT_0_363 : X_AND2 
    port map (
      I0 => UAR1_BYTE_OUT_0_D2_PT_0_0_INV,
      I1 => UAR1_BYTE_OUT_0_FBK,
      O => UAR1_BYTE_OUT_0_D2_PT_0
    );
  UAR1_BYTE_OUT_0_D2_PT_1_364 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_9_FBK,
      O => UAR1_BYTE_OUT_0_D2_PT_1
    );
  UAR1_BYTE_OUT_0_D2_365 : X_OR2 
    port map (
      I0 => UAR1_BYTE_OUT_0_D2_PT_0,
      I1 => UAR1_BYTE_OUT_0_D2_PT_1,
      O => UAR1_BYTE_OUT_0_D2
    );
  UAR1_BYTE_OUT_0_XOR : X_XOR2 
    port map (
      I0 => UAR1_BYTE_OUT_0_D1,
      I1 => UAR1_BYTE_OUT_0_D2,
      O => UAR1_BYTE_OUT_0_D
    );
  UAR1_BYTE_OUT_0_FBK_366 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_0_Q,
      O => UAR1_BYTE_OUT_0_FBK
    );
  CM_PANIC_ON_367 : X_BUF 
    port map (
      I => CM_PANIC_ON_Q,
      O => CM_PANIC_ON
    );
  CM_PANIC_ON_R_OR_PRLD_368 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => CM_PANIC_ON_R_OR_PRLD
    );
  CM_PANIC_ON_REG : X_FF 
    port map (
      I => CM_PANIC_ON_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => CM_PANIC_ON_R_OR_PRLD,
      O => CM_PANIC_ON_Q
    );
  CM_PANIC_ON_D1_369 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => CM_PANIC_ON_D1
    );
  CM_PANIC_ON_D2_PT_0_370 : X_AND2 
    port map (
      I0 => RXD_ACK,
      I1 => RXD_ACK,
      O => CM_PANIC_ON_D2_PT_0
    );
  CM_PANIC_ON_D2_PT_1_371 : X_AND2 
    port map (
      I0 => RXD_2_FBK,
      I1 => RXD_2_FBK,
      O => CM_PANIC_ON_D2_PT_1
    );
  CM_PANIC_ON_D2_PT_2_372 : X_AND2 
    port map (
      I0 => EXP17_EXP,
      I1 => EXP17_EXP,
      O => CM_PANIC_ON_D2_PT_2
    );
  CM_PANIC_ON_D2_PT_3_373 : X_AND2 
    port map (
      I0 => EXP18_EXP,
      I1 => EXP18_EXP,
      O => CM_PANIC_ON_D2_PT_3
    );
  CM_PANIC_ON_D2_PT_4_374 : X_AND2 
    port map (
      I0 => CM_PANIC_ON_D2_PT_4_0_INV,
      I1 => CM_PANIC_ON_D2_PT_4_1_INV,
      O => CM_PANIC_ON_D2_PT_4
    );
  CM_PANIC_ON_D2_PT_5_375 : X_AND2 
    port map (
      I0 => RC_ADDRESS_C(0),
      I1 => CM_PANIC_ON_D2_PT_5_1_INV,
      O => CM_PANIC_ON_D2_PT_5
    );
  CM_PANIC_ON_D2_PT_6_376 : X_AND2 
    port map (
      I0 => CM_PANIC_ON_D2_PT_6_0_INV,
      I1 => RXD_4_FBK,
      O => CM_PANIC_ON_D2_PT_6
    );
  CM_PANIC_ON_D2_377 : X_OR7 
    port map (
      I0 => CM_PANIC_ON_D2_PT_0,
      I1 => CM_PANIC_ON_D2_PT_1,
      I2 => CM_PANIC_ON_D2_PT_2,
      I3 => CM_PANIC_ON_D2_PT_3,
      I4 => CM_PANIC_ON_D2_PT_4,
      I5 => CM_PANIC_ON_D2_PT_5,
      I6 => CM_PANIC_ON_D2_PT_6,
      O => CM_PANIC_ON_D2
    );
  CM_PANIC_ON_D_378 : X_XOR2 
    port map (
      I0 => CM_PANIC_ON_D_TFF,
      I1 => CM_PANIC_ON_Q,
      O => CM_PANIC_ON_D
    );
  CM_PANIC_ON_XOR : X_XOR2 
    port map (
      I0 => CM_PANIC_ON_XOR_0_INV,
      I1 => CM_PANIC_ON_D2,
      O => CM_PANIC_ON_D_TFF
    );
  CM_PANIC_ON_FBK_379 : X_BUF 
    port map (
      I => CM_PANIC_ON_Q,
      O => CM_PANIC_ON_FBK
    );
  EXP17_EXP_PT_0_380 : X_AND2 
    port map (
      I0 => RC_ADDRESS_C(1),
      I1 => EXP17_EXP_PT_0_1_INV,
      O => EXP17_EXP_PT_0
    );
  EXP17_EXP_PT_1_381 : X_AND2 
    port map (
      I0 => EXP17_EXP_PT_1_0_INV,
      I1 => RXD_5_FBK,
      O => EXP17_EXP_PT_1
    );
  EXP17_EXP_PT_2_382 : X_AND2 
    port map (
      I0 => RC_ADDRESS_C(2),
      I1 => EXP17_EXP_PT_2_1_INV,
      O => EXP17_EXP_PT_2
    );
  EXP17_EXP_PT_3_383 : X_AND2 
    port map (
      I0 => EXP17_EXP_PT_3_0_INV,
      I1 => RXD_6_FBK,
      O => EXP17_EXP_PT_3
    );
  EXP17_EXP_PT_4_384 : X_AND2 
    port map (
      I0 => RC_ADDRESS_C(3),
      I1 => EXP17_EXP_PT_4_1_INV,
      O => EXP17_EXP_PT_4
    );
  EXP17_EXP_385 : X_OR5 
    port map (
      I0 => EXP17_EXP_PT_0,
      I1 => EXP17_EXP_PT_1,
      I2 => EXP17_EXP_PT_2,
      I3 => EXP17_EXP_PT_3,
      I4 => EXP17_EXP_PT_4,
      O => EXP17_EXP
    );
  EXP18_EXP_PT_0_386 : X_AND2 
    port map (
      I0 => RXD_0_EXP,
      I1 => RXD_0_EXP,
      O => EXP18_EXP_PT_0
    );
  EXP18_EXP_PT_1_387 : X_AND2 
    port map (
      I0 => RXD_3_FBK,
      I1 => CM_PANIC_ON_FBK,
      O => EXP18_EXP_PT_1
    );
  EXP18_EXP_PT_2_388 : X_AND2 
    port map (
      I0 => EXP18_EXP_PT_2_0_INV,
      I1 => EXP18_EXP_PT_2_1_INV,
      O => EXP18_EXP_PT_2
    );
  EXP18_EXP_PT_3_389 : X_AND2 
    port map (
      I0 => RXD_1_FBK,
      I1 => EXP18_EXP_PT_3_1_INV,
      O => EXP18_EXP_PT_3
    );
  EXP18_EXP_PT_4_390 : X_AND2 
    port map (
      I0 => EXP18_EXP_PT_4_0_INV,
      I1 => RXD_0_FBK,
      O => EXP18_EXP_PT_4
    );
  EXP18_EXP_PT_5_391 : X_AND2 
    port map (
      I0 => EXP18_EXP_PT_5_0_INV,
      I1 => RXD_7_FBK,
      O => EXP18_EXP_PT_5
    );
  EXP18_EXP_392 : X_OR6 
    port map (
      I0 => EXP18_EXP_PT_0,
      I1 => EXP18_EXP_PT_1,
      I2 => EXP18_EXP_PT_2,
      I3 => EXP18_EXP_PT_3,
      I4 => EXP18_EXP_PT_4,
      I5 => EXP18_EXP_PT_5,
      O => EXP18_EXP
    );
  RC_ADDRESS_C_0_Q : X_BUF 
    port map (
      I => RC_ADDRESS(0),
      O => RC_ADDRESS_C(0)
    );
  RXD_4_FBK_393 : X_BUF 
    port map (
      I => RXD_4_Q,
      O => RXD_4_FBK
    );
  RXD_4_R_OR_PRLD_394 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => RXD_4_R_OR_PRLD
    );
  RXD_4_REG : X_FF 
    port map (
      I => RXD_4_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => RXD_4_R_OR_PRLD,
      O => RXD_4_Q
    );
  RXD_4_D1_395 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => RXD_4_D1
    );
  RXD_4_D2_PT_0_396 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_4_D2_PT_0_1_INV,
      I2 => RXD_4_FBK,
      I3 => RXD_4_D2_PT_0_3_INV,
      O => RXD_4_D2_PT_0
    );
  RXD_4_D2_PT_1_397 : X_AND4 
    port map (
      I0 => UAR1_BYTE_AVAIL,
      I1 => RXD_4_D2_PT_1_1_INV,
      I2 => RXD_4_D2_PT_1_2_INV,
      I3 => UAR1_BYTE_OUT(4),
      O => RXD_4_D2_PT_1
    );
  RXD_4_D2_398 : X_OR2 
    port map (
      I0 => RXD_4_D2_PT_0,
      I1 => RXD_4_D2_PT_1,
      O => RXD_4_D2
    );
  RXD_4_D_399 : X_XOR2 
    port map (
      I0 => RXD_4_D_TFF,
      I1 => RXD_4_Q,
      O => RXD_4_D
    );
  RXD_4_XOR : X_XOR2 
    port map (
      I0 => RXD_4_D1,
      I1 => RXD_4_D2,
      O => RXD_4_D_TFF
    );
  UAR1_BYTE_OUT_4_Q_400 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_4_Q,
      O => UAR1_BYTE_OUT(4)
    );
  UAR1_BYTE_OUT_4_R_OR_PRLD_401 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => UAR1_BYTE_OUT_4_R_OR_PRLD
    );
  UAR1_BYTE_OUT_4_REG : X_FF 
    port map (
      I => UAR1_BYTE_OUT_4_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => UAR1_BYTE_OUT_4_R_OR_PRLD,
      O => UAR1_BYTE_OUT_4_Q
    );
  UAR1_BYTE_OUT_4_D1_402 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => UAR1_BYTE_OUT_4_D1
    );
  UAR1_BYTE_OUT_4_D2_PT_0_403 : X_AND2 
    port map (
      I0 => UAR1_BYTE_OUT_4_D2_PT_0_0_INV,
      I1 => UAR1_BYTE_OUT_4_FBK,
      O => UAR1_BYTE_OUT_4_D2_PT_0
    );
  UAR1_BYTE_OUT_4_D2_PT_1_404 : X_AND5 
    port map (
      I0 => UAR1_BIT_DONE,
      I1 => UAR1_BM1_SAMPLED_BITS(0),
      I2 => UAR1_BM1_SAMPLED_BITS(1),
      I3 => UAR1_BM1_SAMPLED_BITS(2),
      I4 => UAR1_BC1_CURRENT_STATE_5_FBK,
      O => UAR1_BYTE_OUT_4_D2_PT_1
    );
  UAR1_BYTE_OUT_4_D2_405 : X_OR2 
    port map (
      I0 => UAR1_BYTE_OUT_4_D2_PT_0,
      I1 => UAR1_BYTE_OUT_4_D2_PT_1,
      O => UAR1_BYTE_OUT_4_D2
    );
  UAR1_BYTE_OUT_4_XOR : X_XOR2 
    port map (
      I0 => UAR1_BYTE_OUT_4_D1,
      I1 => UAR1_BYTE_OUT_4_D2,
      O => UAR1_BYTE_OUT_4_D
    );
  UAR1_BYTE_OUT_4_FBK_406 : X_BUF 
    port map (
      I => UAR1_BYTE_OUT_4_Q,
      O => UAR1_BYTE_OUT_4_FBK
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_Q_407 : X_BUF 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_Q,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0)
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_R_OR_PRLD_408 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_R_OR_PRLD
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_REG : X_FF 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_R_OR_PRLD,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_Q
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D1_409 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D1
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_0_410 : X_AND2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_0
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_1_411 : X_AND2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_1_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_1_1_INV,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_1
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_412 : X_OR2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_0,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_1,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D_413 : X_XOR2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D_TFF,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_Q,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_XOR : X_XOR2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_XOR_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D_TFF
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_414 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_0_INV,
      I1 => LIGHT_VALUE_4_FBK,
      I2 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_2_INV,
      I3 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_3_INV,
      I4 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_4_INV,
      I5 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_5_INV,
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_6_INV,
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_7_INV,
      I8 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_8_INV,
      I9 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_415 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_1_INV,
      I2 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_2_INV,
      I3 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_3_INV,
      I4 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_4_INV,
      I5 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_5_INV,
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_6_INV,
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_7_INV,
      I8 => LIGHT_VALUE(5),
      I9 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_416 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_1_INV,
      I2 => FC1_CNT_3_FBK,
      I3 => FC1_CNT(1),
      I4 => FC1_CNT(2),
      I5 => FC1_CNT_4_FBK,
      I6 => FC1_CNT_5_FBK,
      I7 => FC1_CNT_6_FBK,
      I8 => FC1_CNT(0),
      I9 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_9_INV,
      I10 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_10_INV,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_417 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_1_INV,
      I2 => FC1_CNT_3_FBK,
      I3 => FC1_CNT(1),
      I4 => FC1_CNT(2),
      I5 => FC1_CNT_4_FBK,
      I6 => FC1_CNT_5_FBK,
      I7 => FC1_CNT_6_FBK,
      I8 => FC1_CNT(0),
      I9 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_9_INV,
      I10 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_10_INV,
      I11 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_11_INV,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_418 : X_OR4 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1,
      I2 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2,
      I3 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK_419 : X_BUF 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_Q,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK
    );
  FC1_CNT_3_Q_420 : X_BUF 
    port map (
      I => FC1_CNT_3_Q,
      O => FC1_CNT(3)
    );
  FC1_CNT_3_R_OR_PRLD_421 : X_OR2 
    port map (
      I0 => FC1_CNT_3_RSTF,
      I1 => PRLD,
      O => FC1_CNT_3_R_OR_PRLD
    );
  FC1_CNT_3_REG : X_FF 
    port map (
      I => FC1_CNT_3_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => FC1_CNT_3_R_OR_PRLD,
      O => FC1_CNT_3_Q
    );
  FC1_CNT_3_RSTF_PT_0_422 : X_AND2 
    port map (
      I0 => FC1_CNT_3_RSTF_PT_0_0_INV,
      I1 => FC1_CNT_3_RSTF_PT_0_1_INV,
      O => FC1_CNT_3_RSTF_PT_0
    );
  FC1_CNT_3_RSTF_423 : X_OR2 
    port map (
      I0 => FC1_CNT_3_RSTF_PT_0,
      I1 => FC1_CNT_3_RSTF_PT_0,
      O => FC1_CNT_3_RSTF
    );
  FC1_CNT_3_D1_424 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => FC1_CNT_3_D1
    );
  FC1_CNT_3_D2_PT_0_425 : X_AND2 
    port map (
      I0 => EXP4_EXP,
      I1 => EXP4_EXP,
      O => FC1_CNT_3_D2_PT_0
    );
  FC1_CNT_3_D2_PT_1_426 : X_AND4 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => LIGHT_VALUE(5),
      I2 => LIGHT_VALUE(3),
      I3 => LIGHT_VALUE(2),
      O => FC1_CNT_3_D2_PT_1
    );
  FC1_CNT_3_D2_PT_2_427 : X_AND16 
    port map (
      I0 => FC1_CNT_3_D2_PT_2_0_INV,
      I1 => FC1_CNT_3_D2_PT_2_1_INV,
      I2 => FC1_CNT_3_D2_PT_2_2_INV,
      I3 => FC1_CNT_3_D2_PT_2_3_INV,
      I4 => FC1_CNT_3_D2_PT_2_4_INV,
      I5 => FC1_CNT_3_D2_PT_2_5_INV,
      I6 => FC1_CNT_3_D2_PT_2_6_INV,
      I7 => FC1_CNT_3_D2_PT_2_7_INV,
      I8 => FC1_CNT_3_D2_PT_2_8_INV,
      I9 => FC1_CNT_3_D2_PT_2_9_INV,
      I10 => FC1_CNT_3_D2_PT_2_10_INV,
      I11 => FC1_CNT_3_D2_PT_2_11_INV,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_3_D2_PT_2
    );
  FC1_CNT_3_D2_428 : X_OR3 
    port map (
      I0 => FC1_CNT_3_D2_PT_0,
      I1 => FC1_CNT_3_D2_PT_1,
      I2 => FC1_CNT_3_D2_PT_2,
      O => FC1_CNT_3_D2
    );
  FC1_CNT_3_D_429 : X_XOR2 
    port map (
      I0 => FC1_CNT_3_D_TFF,
      I1 => FC1_CNT_3_Q,
      O => FC1_CNT_3_D
    );
  FC1_CNT_3_XOR : X_XOR2 
    port map (
      I0 => FC1_CNT_3_XOR_0_INV,
      I1 => FC1_CNT_3_D2,
      O => FC1_CNT_3_D_TFF
    );
  FC1_CNT_3_EXP_PT_0_430 : X_AND16 
    port map (
      I0 => FC1_CNT_3_EXP_PT_0_0_INV,
      I1 => FC1_CNT_3_EXP_PT_0_1_INV,
      I2 => FC1_CNT_3_EXP_PT_0_2_INV,
      I3 => FC1_CNT_3_EXP_PT_0_3_INV,
      I4 => FC1_CNT_3_EXP_PT_0_4_INV,
      I5 => FC1_CNT_3_EXP_PT_0_5_INV,
      I6 => FC1_CNT_3_EXP_PT_0_6_INV,
      I7 => LIGHT_VALUE(3),
      I8 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I9 => VCC,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_3_EXP_PT_0
    );
  FC1_CNT_3_EXP_PT_1_431 : X_AND16 
    port map (
      I0 => FC1_CNT_3_EXP_PT_1_0_INV,
      I1 => FC1_CNT_3_EXP_PT_1_1_INV,
      I2 => FC1_CNT_3_EXP_PT_1_2_INV,
      I3 => FC1_CNT_3_EXP_PT_1_3_INV,
      I4 => FC1_CNT_3_EXP_PT_1_4_INV,
      I5 => FC1_CNT_3_EXP_PT_1_5_INV,
      I6 => FC1_CNT_3_EXP_PT_1_6_INV,
      I7 => LIGHT_VALUE(1),
      I8 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I9 => VCC,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_3_EXP_PT_1
    );
  FC1_CNT_3_EXP_432 : X_OR2 
    port map (
      I0 => FC1_CNT_3_EXP_PT_0,
      I1 => FC1_CNT_3_EXP_PT_1,
      O => FC1_CNT_3_EXP
    );
  FC1_CNT_3_FBK_433 : X_BUF 
    port map (
      I => FC1_CNT_3_Q,
      O => FC1_CNT_3_FBK
    );
  EXP4_EXP_PT_0_434 : X_AND2 
    port map (
      I0 => FC1_CNT_7_EXP,
      I1 => FC1_CNT_7_EXP,
      O => EXP4_EXP_PT_0
    );
  EXP4_EXP_PT_1_435 : X_AND2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP4_EXP_PT_1
    );
  EXP4_EXP_PT_2_436 : X_AND2 
    port map (
      I0 => EXP4_EXP_PT_2_0_INV,
      I1 => FC1_CNT(0),
      O => EXP4_EXP_PT_2
    );
  EXP4_EXP_PT_3_437 : X_AND2 
    port map (
      I0 => FC1_CNT(1),
      I1 => EXP4_EXP_PT_3_1_INV,
      O => EXP4_EXP_PT_3
    );
  EXP4_EXP_PT_4_438 : X_AND3 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => LIGHT_VALUE_4_FBK,
      I2 => LIGHT_VALUE(5),
      O => EXP4_EXP_PT_4
    );
  EXP4_EXP_PT_5_439 : X_AND4 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => LIGHT_VALUE(5),
      I2 => LIGHT_VALUE(3),
      I3 => LIGHT_VALUE(1),
      O => EXP4_EXP_PT_5
    );
  EXP4_EXP_440 : X_OR6 
    port map (
      I0 => EXP4_EXP_PT_0,
      I1 => EXP4_EXP_PT_1,
      I2 => EXP4_EXP_PT_2,
      I3 => EXP4_EXP_PT_3,
      I4 => EXP4_EXP_PT_4,
      I5 => EXP4_EXP_PT_5,
      O => EXP4_EXP
    );
  FC1_CNT_7_Q_441 : X_BUF 
    port map (
      I => FC1_CNT_7_Q,
      O => FC1_CNT(7)
    );
  FC1_CNT_7_R_OR_PRLD_442 : X_OR2 
    port map (
      I0 => FC1_CNT_7_RSTF,
      I1 => PRLD,
      O => FC1_CNT_7_R_OR_PRLD
    );
  FC1_CNT_7_REG : X_FF 
    port map (
      I => FC1_CNT_7_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => FC1_CNT_7_R_OR_PRLD,
      O => FC1_CNT_7_Q
    );
  FC1_CNT_7_RSTF_PT_0_443 : X_AND2 
    port map (
      I0 => FC1_CNT_7_RSTF_PT_0_0_INV,
      I1 => FC1_CNT_7_RSTF_PT_0_1_INV,
      O => FC1_CNT_7_RSTF_PT_0
    );
  FC1_CNT_7_RSTF_444 : X_OR2 
    port map (
      I0 => FC1_CNT_7_RSTF_PT_0,
      I1 => FC1_CNT_7_RSTF_PT_0,
      O => FC1_CNT_7_RSTF
    );
  FC1_CNT_7_D1_445 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => FC1_CNT_7_D1
    );
  FC1_CNT_7_D2_PT_0_446 : X_AND2 
    port map (
      I0 => EXP3_EXP,
      I1 => EXP3_EXP,
      O => FC1_CNT_7_D2_PT_0
    );
  FC1_CNT_7_D2_PT_1_447 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => FC1_CNT_3_FBK,
      I2 => FC1_CNT(1),
      I3 => FC1_CNT(2),
      I4 => FC1_CNT_4_FBK,
      I5 => FC1_CNT_5_FBK,
      I6 => FC1_CNT_6_FBK,
      I7 => FC1_CNT(0),
      I8 => FC1_CNT_7_D2_PT_1_8_INV,
      I9 => FC1_CNT_7_D2_PT_1_9_INV,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_7_D2_PT_1
    );
  FC1_CNT_7_D2_448 : X_OR2 
    port map (
      I0 => FC1_CNT_7_D2_PT_0,
      I1 => FC1_CNT_7_D2_PT_1,
      O => FC1_CNT_7_D2
    );
  FC1_CNT_7_D_449 : X_XOR2 
    port map (
      I0 => FC1_CNT_7_D_TFF,
      I1 => FC1_CNT_7_Q,
      O => FC1_CNT_7_D
    );
  FC1_CNT_7_XOR : X_XOR2 
    port map (
      I0 => FC1_CNT_7_D1,
      I1 => FC1_CNT_7_D2,
      O => FC1_CNT_7_D_TFF
    );
  FC1_CNT_7_EXP_PT_0_450 : X_AND2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => FC1_CNT_7_EXP_PT_0_1_INV,
      O => FC1_CNT_7_EXP_PT_0
    );
  FC1_CNT_7_EXP_PT_1_451 : X_AND2 
    port map (
      I0 => FC1_CNT_7_EXP_PT_1_0_INV,
      I1 => FC1_CNT_7_EXP_PT_1_1_INV,
      O => FC1_CNT_7_EXP_PT_1
    );
  FC1_CNT_7_EXP_PT_2_452 : X_AND2 
    port map (
      I0 => FC1_CNT_7_EXP_PT_2_0_INV,
      I1 => FC1_CNT(2),
      O => FC1_CNT_7_EXP_PT_2
    );
  FC1_CNT_7_EXP_453 : X_OR3 
    port map (
      I0 => FC1_CNT_7_EXP_PT_0,
      I1 => FC1_CNT_7_EXP_PT_1,
      I2 => FC1_CNT_7_EXP_PT_2,
      O => FC1_CNT_7_EXP
    );
  FC1_CNT_7_FBK_454 : X_BUF 
    port map (
      I => FC1_CNT_7_Q,
      O => FC1_CNT_7_FBK
    );
  EXP3_EXP_PT_0_455 : X_AND2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP,
      O => EXP3_EXP_PT_0
    );
  EXP3_EXP_PT_1_456 : X_AND16 
    port map (
      I0 => EXP3_EXP_PT_1_0_INV,
      I1 => EXP3_EXP_PT_1_1_INV,
      I2 => EXP3_EXP_PT_1_2_INV,
      I3 => EXP3_EXP_PT_1_3_INV,
      I4 => EXP3_EXP_PT_1_4_INV,
      I5 => EXP3_EXP_PT_1_5_INV,
      I6 => EXP3_EXP_PT_1_6_INV,
      I7 => EXP3_EXP_PT_1_7_INV,
      I8 => LIGHT_VALUE(3),
      I9 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP3_EXP_PT_1
    );
  EXP3_EXP_PT_2_457 : X_AND16 
    port map (
      I0 => EXP3_EXP_PT_2_0_INV,
      I1 => EXP3_EXP_PT_2_1_INV,
      I2 => EXP3_EXP_PT_2_2_INV,
      I3 => EXP3_EXP_PT_2_3_INV,
      I4 => EXP3_EXP_PT_2_4_INV,
      I5 => EXP3_EXP_PT_2_5_INV,
      I6 => EXP3_EXP_PT_2_6_INV,
      I7 => EXP3_EXP_PT_2_7_INV,
      I8 => LIGHT_VALUE(1),
      I9 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP3_EXP_PT_2
    );
  EXP3_EXP_PT_3_458 : X_AND16 
    port map (
      I0 => EXP3_EXP_PT_3_0_INV,
      I1 => EXP3_EXP_PT_3_1_INV,
      I2 => EXP3_EXP_PT_3_2_INV,
      I3 => EXP3_EXP_PT_3_3_INV,
      I4 => EXP3_EXP_PT_3_4_INV,
      I5 => EXP3_EXP_PT_3_5_INV,
      I6 => EXP3_EXP_PT_3_6_INV,
      I7 => EXP3_EXP_PT_3_7_INV,
      I8 => LIGHT_VALUE(2),
      I9 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP3_EXP_PT_3
    );
  EXP3_EXP_PT_4_459 : X_AND16 
    port map (
      I0 => EXP3_EXP_PT_4_0_INV,
      I1 => EXP3_EXP_PT_4_1_INV,
      I2 => EXP3_EXP_PT_4_2_INV,
      I3 => EXP3_EXP_PT_4_3_INV,
      I4 => EXP3_EXP_PT_4_4_INV,
      I5 => EXP3_EXP_PT_4_5_INV,
      I6 => EXP3_EXP_PT_4_6_INV,
      I7 => EXP3_EXP_PT_4_7_INV,
      I8 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I9 => LIGHT_VALUE(0),
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP3_EXP_PT_4
    );
  EXP3_EXP_PT_5_460 : X_AND16 
    port map (
      I0 => EXP3_EXP_PT_5_0_INV,
      I1 => EXP3_EXP_PT_5_1_INV,
      I2 => EXP3_EXP_PT_5_2_INV,
      I3 => EXP3_EXP_PT_5_3_INV,
      I4 => EXP3_EXP_PT_5_4_INV,
      I5 => EXP3_EXP_PT_5_5_INV,
      I6 => EXP3_EXP_PT_5_6_INV,
      I7 => EXP3_EXP_PT_5_7_INV,
      I8 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I9 => FC1_CNT_7_FBK,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP3_EXP_PT_5
    );
  EXP3_EXP_461 : X_OR6 
    port map (
      I0 => EXP3_EXP_PT_0,
      I1 => EXP3_EXP_PT_1,
      I2 => EXP3_EXP_PT_2,
      I3 => EXP3_EXP_PT_3,
      I4 => EXP3_EXP_PT_4,
      I5 => EXP3_EXP_PT_5,
      O => EXP3_EXP
    );
  FC1_CNT_1_Q_462 : X_BUF 
    port map (
      I => FC1_CNT_1_Q,
      O => FC1_CNT(1)
    );
  FC1_CNT_1_R_OR_PRLD_463 : X_OR2 
    port map (
      I0 => FC1_CNT_1_RSTF,
      I1 => PRLD,
      O => FC1_CNT_1_R_OR_PRLD
    );
  FC1_CNT_1_REG : X_FF 
    port map (
      I => FC1_CNT_1_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => FC1_CNT_1_R_OR_PRLD,
      O => FC1_CNT_1_Q
    );
  FC1_CNT_1_RSTF_PT_0_464 : X_AND2 
    port map (
      I0 => FC1_CNT_1_RSTF_PT_0_0_INV,
      I1 => FC1_CNT_1_RSTF_PT_0_1_INV,
      O => FC1_CNT_1_RSTF_PT_0
    );
  FC1_CNT_1_RSTF_465 : X_OR2 
    port map (
      I0 => FC1_CNT_1_RSTF_PT_0,
      I1 => FC1_CNT_1_RSTF_PT_0,
      O => FC1_CNT_1_RSTF
    );
  FC1_CNT_1_D1_466 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => FC1_CNT_1_D1
    );
  FC1_CNT_1_D2_PT_0_467 : X_AND2 
    port map (
      I0 => FC1_CNT_0_EXP,
      I1 => FC1_CNT_0_EXP,
      O => FC1_CNT_1_D2_PT_0
    );
  FC1_CNT_1_D2_PT_1_468 : X_AND3 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I1 => LIGHT_VALUE_5_FBK,
      I2 => LIGHT_VALUE(4),
      O => FC1_CNT_1_D2_PT_1
    );
  FC1_CNT_1_D2_PT_2_469 : X_AND4 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I1 => LIGHT_VALUE_5_FBK,
      I2 => LIGHT_VALUE_1_FBK,
      I3 => LIGHT_VALUE_3_FBK,
      O => FC1_CNT_1_D2_PT_2
    );
  FC1_CNT_1_D2_PT_3_470 : X_AND4 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I1 => LIGHT_VALUE_5_FBK,
      I2 => LIGHT_VALUE_2_FBK,
      I3 => LIGHT_VALUE_3_FBK,
      O => FC1_CNT_1_D2_PT_3
    );
  FC1_CNT_1_D2_PT_4_471 : X_AND16 
    port map (
      I0 => FC1_CNT_1_D2_PT_4_0_INV,
      I1 => FC1_CNT_1_D2_PT_4_1_INV,
      I2 => FC1_CNT_1_D2_PT_4_2_INV,
      I3 => FC1_CNT_1_D2_PT_4_3_INV,
      I4 => FC1_CNT_1_D2_PT_4_4_INV,
      I5 => FC1_CNT_1_D2_PT_4_5_INV,
      I6 => FC1_CNT_1_D2_PT_4_6_INV,
      I7 => FC1_CNT_1_D2_PT_4_7_INV,
      I8 => FC1_CNT_1_D2_PT_4_8_INV,
      I9 => FC1_CNT_1_D2_PT_4_9_INV,
      I10 => FC1_CNT_1_D2_PT_4_10_INV,
      I11 => FC1_CNT_1_D2_PT_4_11_INV,
      I12 => FC1_CNT_1_D2_PT_4_12_INV,
      I13 => FC1_CNT_1_D2_PT_4_13_INV,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_1_D2_PT_4
    );
  FC1_CNT_1_D2_472 : X_OR5 
    port map (
      I0 => FC1_CNT_1_D2_PT_0,
      I1 => FC1_CNT_1_D2_PT_1,
      I2 => FC1_CNT_1_D2_PT_2,
      I3 => FC1_CNT_1_D2_PT_3,
      I4 => FC1_CNT_1_D2_PT_4,
      O => FC1_CNT_1_D2
    );
  FC1_CNT_1_D_473 : X_XOR2 
    port map (
      I0 => FC1_CNT_1_D_TFF,
      I1 => FC1_CNT_1_Q,
      O => FC1_CNT_1_D
    );
  FC1_CNT_1_XOR : X_XOR2 
    port map (
      I0 => FC1_CNT_1_XOR_0_INV,
      I1 => FC1_CNT_1_D2,
      O => FC1_CNT_1_D_TFF
    );
  FC1_CNT_1_FBK_474 : X_BUF 
    port map (
      I => FC1_CNT_1_Q,
      O => FC1_CNT_1_FBK
    );
  FC1_CNT_0_Q_475 : X_BUF 
    port map (
      I => FC1_CNT_0_Q,
      O => FC1_CNT(0)
    );
  FC1_CNT_0_R_OR_PRLD_476 : X_OR2 
    port map (
      I0 => FC1_CNT_0_RSTF,
      I1 => PRLD,
      O => FC1_CNT_0_R_OR_PRLD
    );
  FC1_CNT_0_REG : X_FF 
    port map (
      I => FC1_CNT_0_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => FC1_CNT_0_R_OR_PRLD,
      O => FC1_CNT_0_Q
    );
  FC1_CNT_0_RSTF_PT_0_477 : X_AND2 
    port map (
      I0 => FC1_CNT_0_RSTF_PT_0_0_INV,
      I1 => FC1_CNT_0_RSTF_PT_0_1_INV,
      O => FC1_CNT_0_RSTF_PT_0
    );
  FC1_CNT_0_RSTF_478 : X_OR2 
    port map (
      I0 => FC1_CNT_0_RSTF_PT_0,
      I1 => FC1_CNT_0_RSTF_PT_0,
      O => FC1_CNT_0_RSTF
    );
  FC1_CNT_0_D1_479 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => FC1_CNT_0_D1
    );
  FC1_CNT_0_D2_PT_0_480 : X_AND2 
    port map (
      I0 => EXP12_EXP,
      I1 => EXP12_EXP,
      O => FC1_CNT_0_D2_PT_0
    );
  FC1_CNT_0_D2_PT_1_481 : X_AND2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => FC1_CNT_0_D2_PT_1
    );
  FC1_CNT_0_D2_482 : X_OR2 
    port map (
      I0 => FC1_CNT_0_D2_PT_0,
      I1 => FC1_CNT_0_D2_PT_1,
      O => FC1_CNT_0_D2
    );
  FC1_CNT_0_D_483 : X_XOR2 
    port map (
      I0 => FC1_CNT_0_D_TFF,
      I1 => FC1_CNT_0_Q,
      O => FC1_CNT_0_D
    );
  FC1_CNT_0_XOR : X_XOR2 
    port map (
      I0 => FC1_CNT_0_XOR_0_INV,
      I1 => FC1_CNT_0_D2,
      O => FC1_CNT_0_D_TFF
    );
  FC1_CNT_0_EXP_PT_0_484 : X_AND2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => FC1_CNT_0_EXP_PT_0
    );
  FC1_CNT_0_EXP_PT_1_485 : X_AND2 
    port map (
      I0 => FC1_CNT_0_EXP_PT_1_0_INV,
      I1 => FC1_CNT_0_EXP_PT_1_1_INV,
      O => FC1_CNT_0_EXP_PT_1
    );
  FC1_CNT_0_EXP_PT_2_486 : X_AND2 
    port map (
      I0 => FC1_CNT_0_EXP_PT_2_0_INV,
      I1 => FC1_CNT_0_FBK,
      O => FC1_CNT_0_EXP_PT_2
    );
  FC1_CNT_0_EXP_487 : X_OR3 
    port map (
      I0 => FC1_CNT_0_EXP_PT_0,
      I1 => FC1_CNT_0_EXP_PT_1,
      I2 => FC1_CNT_0_EXP_PT_2,
      O => FC1_CNT_0_EXP
    );
  FC1_CNT_0_FBK_488 : X_BUF 
    port map (
      I => FC1_CNT_0_Q,
      O => FC1_CNT_0_FBK
    );
  EXP12_EXP_PT_0_489 : X_AND2 
    port map (
      I0 => EXP12_EXP_PT_0_0_INV,
      I1 => EXP12_EXP_PT_0_1_INV,
      O => EXP12_EXP_PT_0
    );
  EXP12_EXP_PT_1_490 : X_AND3 
    port map (
      I0 => EXP12_EXP_PT_1_0_INV,
      I1 => LIGHT_VALUE_5_FBK,
      I2 => LIGHT_VALUE(4),
      O => EXP12_EXP_PT_1
    );
  EXP12_EXP_PT_2_491 : X_AND4 
    port map (
      I0 => EXP12_EXP_PT_2_0_INV,
      I1 => LIGHT_VALUE_5_FBK,
      I2 => LIGHT_VALUE_1_FBK,
      I3 => LIGHT_VALUE_3_FBK,
      O => EXP12_EXP_PT_2
    );
  EXP12_EXP_PT_3_492 : X_AND4 
    port map (
      I0 => EXP12_EXP_PT_3_0_INV,
      I1 => LIGHT_VALUE_5_FBK,
      I2 => LIGHT_VALUE_2_FBK,
      I3 => LIGHT_VALUE_3_FBK,
      O => EXP12_EXP_PT_3
    );
  EXP12_EXP_PT_4_493 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => EXP12_EXP_PT_4_1_INV,
      I2 => EXP12_EXP_PT_4_2_INV,
      I3 => EXP12_EXP_PT_4_3_INV,
      I4 => EXP12_EXP_PT_4_4_INV,
      I5 => EXP12_EXP_PT_4_5_INV,
      I6 => EXP12_EXP_PT_4_6_INV,
      I7 => EXP12_EXP_PT_4_7_INV,
      I8 => EXP12_EXP_PT_4_8_INV,
      I9 => EXP12_EXP_PT_4_9_INV,
      I10 => EXP12_EXP_PT_4_10_INV,
      I11 => EXP12_EXP_PT_4_11_INV,
      I12 => EXP12_EXP_PT_4_12_INV,
      I13 => EXP12_EXP_PT_4_13_INV,
      I14 => EXP12_EXP_PT_4_14_INV,
      I15 => VCC,
      O => EXP12_EXP_PT_4
    );
  EXP12_EXP_494 : X_OR5 
    port map (
      I0 => EXP12_EXP_PT_0,
      I1 => EXP12_EXP_PT_1,
      I2 => EXP12_EXP_PT_2,
      I3 => EXP12_EXP_PT_3,
      I4 => EXP12_EXP_PT_4,
      O => EXP12_EXP
    );
  LIGHT_VALUE_5_Q_495 : X_BUF 
    port map (
      I => LIGHT_VALUE_5_Q,
      O => LIGHT_VALUE(5)
    );
  LIGHT_VALUE_5_REG : X_FF 
    port map (
      I => LIGHT_VALUE_5_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => LIGHT_VALUE_5_SETF,
      RST => PRLD,
      O => LIGHT_VALUE_5_Q
    );
  LIGHT_VALUE_5_SETF_PT_0_496 : X_AND2 
    port map (
      I0 => LIGHT_VALUE_5_SETF_PT_0_0_INV,
      I1 => LIGHT_VALUE_5_SETF_PT_0_1_INV,
      O => LIGHT_VALUE_5_SETF_PT_0
    );
  LIGHT_VALUE_5_SETF_497 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_5_SETF_PT_0,
      I1 => LIGHT_VALUE_5_SETF_PT_0,
      O => LIGHT_VALUE_5_SETF
    );
  LIGHT_VALUE_5_D1_498 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => LIGHT_VALUE_5_D1
    );
  LIGHT_VALUE_5_D2_PT_0_499 : X_AND2 
    port map (
      I0 => TD1_CNT_0_EXP,
      I1 => TD1_CNT_0_EXP,
      O => LIGHT_VALUE_5_D2_PT_0
    );
  LIGHT_VALUE_5_D2_PT_1_500 : X_AND16 
    port map (
      I0 => LIGHT_VALUE_5_D2_PT_1_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I2 => LIGHT_VALUE_5_D2_PT_1_2_INV,
      I3 => FC1_CNT_1_FBK,
      I4 => FC1_CNT_2_FBK,
      I5 => FC1_CNT_0_FBK,
      I6 => FC1_CNT(3),
      I7 => FC1_CNT(4),
      I8 => FC1_CNT(5),
      I9 => FC1_CNT(6),
      I10 => FC1_CNT(7),
      I11 => LIGHT_VALUE_1_FBK,
      I12 => LIGHT_VALUE_2_FBK,
      I13 => LIGHT_VALUE_0_FBK,
      I14 => LIGHT_VALUE_3_FBK,
      I15 => LIGHT_VALUE(4),
      O => LIGHT_VALUE_5_D2_PT_1
    );
  LIGHT_VALUE_5_D2_501 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_5_D2_PT_0,
      I1 => LIGHT_VALUE_5_D2_PT_1,
      O => LIGHT_VALUE_5_D2
    );
  LIGHT_VALUE_5_D_502 : X_XOR2 
    port map (
      I0 => LIGHT_VALUE_5_D_TFF,
      I1 => LIGHT_VALUE_5_Q,
      O => LIGHT_VALUE_5_D
    );
  LIGHT_VALUE_5_XOR : X_XOR2 
    port map (
      I0 => LIGHT_VALUE_5_D1,
      I1 => LIGHT_VALUE_5_D2,
      O => LIGHT_VALUE_5_D_TFF
    );
  LIGHT_VALUE_5_EXP_PT_0_503 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => LIGHT_VALUE_5_EXP_PT_0_1_INV,
      I2 => LIGHT_VALUE_5_FBK,
      I3 => LIGHT_VALUE_5_EXP_PT_0_3_INV,
      I4 => LIGHT_VALUE_5_EXP_PT_0_4_INV,
      I5 => LIGHT_VALUE_5_EXP_PT_0_5_INV,
      I6 => LIGHT_VALUE_5_EXP_PT_0_6_INV,
      I7 => LIGHT_VALUE_5_EXP_PT_0_7_INV,
      I8 => LIGHT_VALUE_5_EXP_PT_0_8_INV,
      I9 => LIGHT_VALUE_5_EXP_PT_0_9_INV,
      I10 => LIGHT_VALUE_5_EXP_PT_0_10_INV,
      I11 => LIGHT_VALUE_5_EXP_PT_0_11_INV,
      I12 => LIGHT_VALUE_5_EXP_PT_0_12_INV,
      I13 => LIGHT_VALUE_5_EXP_PT_0_13_INV,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_5_EXP_PT_0
    );
  LIGHT_VALUE_5_EXP_PT_1_504 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => LIGHT_VALUE_5_EXP_PT_1_1_INV,
      I2 => LIGHT_VALUE_5_EXP_PT_1_2_INV,
      I3 => LIGHT_VALUE_5_EXP_PT_1_3_INV,
      I4 => LIGHT_VALUE_5_EXP_PT_1_4_INV,
      I5 => LIGHT_VALUE_5_EXP_PT_1_5_INV,
      I6 => LIGHT_VALUE_5_EXP_PT_1_6_INV,
      I7 => LIGHT_VALUE_5_EXP_PT_1_7_INV,
      I8 => LIGHT_VALUE_5_EXP_PT_1_8_INV,
      I9 => LIGHT_VALUE_5_EXP_PT_1_9_INV,
      I10 => LIGHT_VALUE_5_EXP_PT_1_10_INV,
      I11 => LIGHT_VALUE_5_EXP_PT_1_11_INV,
      I12 => LIGHT_VALUE_5_EXP_PT_1_12_INV,
      I13 => LIGHT_VALUE(4),
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_5_EXP_PT_1
    );
  LIGHT_VALUE_5_EXP_PT_2_505 : X_AND16 
    port map (
      I0 => LIGHT_VALUE_5_EXP_PT_2_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I2 => FC1_CNT_1_FBK,
      I3 => FC1_CNT_2_FBK,
      I4 => FC1_CNT_0_FBK,
      I5 => FC1_CNT(3),
      I6 => FC1_CNT(4),
      I7 => FC1_CNT(5),
      I8 => FC1_CNT(6),
      I9 => FC1_CNT(7),
      I10 => LIGHT_VALUE_1_FBK,
      I11 => LIGHT_VALUE_2_FBK,
      I12 => LIGHT_VALUE_0_FBK,
      I13 => LIGHT_VALUE_5_EXP_PT_2_13_INV,
      I14 => LIGHT_VALUE_5_EXP_PT_2_14_INV,
      I15 => VCC,
      O => LIGHT_VALUE_5_EXP_PT_2
    );
  LIGHT_VALUE_5_EXP_506 : X_OR3 
    port map (
      I0 => LIGHT_VALUE_5_EXP_PT_0,
      I1 => LIGHT_VALUE_5_EXP_PT_1,
      I2 => LIGHT_VALUE_5_EXP_PT_2,
      O => LIGHT_VALUE_5_EXP
    );
  LIGHT_VALUE_5_FBK_507 : X_BUF 
    port map (
      I => LIGHT_VALUE_5_Q,
      O => LIGHT_VALUE_5_FBK
    );
  TD1_CNT_0_Q_508 : X_BUF 
    port map (
      I => TD1_CNT_0_Q,
      O => TD1_CNT_0_Q_2
    );
  TD1_CNT_0_R_OR_PRLD_509 : X_OR2 
    port map (
      I0 => TD1_CNT_0_RSTF,
      I1 => PRLD,
      O => TD1_CNT_0_R_OR_PRLD
    );
  TD1_CNT_0_REG : X_FF 
    port map (
      I => TD1_CNT_0_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => TD1_CNT_0_R_OR_PRLD,
      O => TD1_CNT_0_Q
    );
  TD1_CNT_0_RSTF_PT_0_510 : X_AND2 
    port map (
      I0 => TD1_CNT_0_RSTF_PT_0_0_INV,
      I1 => TD1_CNT_0_RSTF_PT_0_1_INV,
      O => TD1_CNT_0_RSTF_PT_0
    );
  TD1_CNT_0_RSTF_511 : X_OR2 
    port map (
      I0 => TD1_CNT_0_RSTF_PT_0,
      I1 => TD1_CNT_0_RSTF_PT_0,
      O => TD1_CNT_0_RSTF
    );
  TD1_CNT_0_D1_512 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => TD1_CNT_0_D1
    );
  TD1_CNT_0_D2_PT_0_513 : X_AND2 
    port map (
      I0 => TD1_CNT_0_D2_PT_0_0_INV,
      I1 => TD1_CNT_0_D2_PT_0_1_INV,
      O => TD1_CNT_0_D2_PT_0
    );
  TD1_CNT_0_D2_514 : X_OR2 
    port map (
      I0 => TD1_CNT_0_D2_PT_0,
      I1 => TD1_CNT_0_D2_PT_0,
      O => TD1_CNT_0_D2
    );
  TD1_CNT_0_XOR : X_XOR2 
    port map (
      I0 => TD1_CNT_0_D1,
      I1 => TD1_CNT_0_D2,
      O => TD1_CNT_0_D
    );
  TD1_CNT_0_EXP_PT_0_515 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => TD1_CNT_0_EXP_PT_0_1_INV,
      I2 => LIGHT_VALUE_5_FBK,
      I3 => TD1_CNT_0_EXP_PT_0_3_INV,
      I4 => TD1_CNT_0_EXP_PT_0_4_INV,
      I5 => TD1_CNT_0_EXP_PT_0_5_INV,
      I6 => TD1_CNT_0_EXP_PT_0_6_INV,
      I7 => TD1_CNT_0_EXP_PT_0_7_INV,
      I8 => TD1_CNT_0_EXP_PT_0_8_INV,
      I9 => TD1_CNT_0_EXP_PT_0_9_INV,
      I10 => TD1_CNT_0_EXP_PT_0_10_INV,
      I11 => TD1_CNT_0_EXP_PT_0_11_INV,
      I12 => TD1_CNT_0_EXP_PT_0_12_INV,
      I13 => TD1_CNT_0_EXP_PT_0_13_INV,
      I14 => TD1_CNT_0_EXP_PT_0_14_INV,
      I15 => TD1_CNT_0_EXP_PT_0_15_INV,
      O => TD1_CNT_0_EXP_PT_0
    );
  TD1_CNT_0_EXP_516 : X_OR2 
    port map (
      I0 => TD1_CNT_0_EXP_PT_0,
      I1 => TD1_CNT_0_EXP_PT_0,
      O => TD1_CNT_0_EXP
    );
  TD1_CNT_0_FBK_517 : X_BUF 
    port map (
      I => TD1_CNT_0_Q,
      O => TD1_CNT_0_FBK
    );
  TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM_518 : X_BUF 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_Q,
      O => TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM
    );
  TD1_CNT_5_TD1_CNT_5_SETF_INT_REG : X_BUF 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_D,
      O => TD1_CNT_5_TD1_CNT_5_SETF_INT_Q
    );
  TD1_CNT_5_TD1_CNT_5_SETF_INT_D1_519 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => TD1_CNT_5_TD1_CNT_5_SETF_INT_D1
    );
  TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0_520 : X_AND2 
    port map (
      I0 => TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0_0_INV,
      I1 => TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0_1_INV,
      O => TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0
    );
  TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_521 : X_OR2 
    port map (
      I0 => TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0,
      I1 => TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0,
      O => TD1_CNT_5_TD1_CNT_5_SETF_INT_D2
    );
  TD1_CNT_5_TD1_CNT_5_SETF_INT_XOR : X_XOR2 
    port map (
      I0 => TD1_CNT_5_TD1_CNT_5_SETF_INT_D1,
      I1 => TD1_CNT_5_TD1_CNT_5_SETF_INT_D2,
      O => TD1_CNT_5_TD1_CNT_5_SETF_INT_D
    );
  TD1_CNT_5_TD1_CNT_5_SETF_INT_FBK_522 : X_BUF 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_Q,
      O => TD1_CNT_5_TD1_CNT_5_SETF_INT_FBK
    );
  ZERO_DETECT_C_523 : X_BUF 
    port map (
      I => ZERO_DETECT,
      O => ZERO_DETECT_C
    );
  FC1_CNT_2_Q_524 : X_BUF 
    port map (
      I => FC1_CNT_2_Q,
      O => FC1_CNT(2)
    );
  FC1_CNT_2_R_OR_PRLD_525 : X_OR2 
    port map (
      I0 => FC1_CNT_2_RSTF,
      I1 => PRLD,
      O => FC1_CNT_2_R_OR_PRLD
    );
  FC1_CNT_2_REG : X_FF 
    port map (
      I => FC1_CNT_2_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => FC1_CNT_2_R_OR_PRLD,
      O => FC1_CNT_2_Q
    );
  FC1_CNT_2_RSTF_PT_0_526 : X_AND2 
    port map (
      I0 => FC1_CNT_2_RSTF_PT_0_0_INV,
      I1 => FC1_CNT_2_RSTF_PT_0_1_INV,
      O => FC1_CNT_2_RSTF_PT_0
    );
  FC1_CNT_2_RSTF_527 : X_OR2 
    port map (
      I0 => FC1_CNT_2_RSTF_PT_0,
      I1 => FC1_CNT_2_RSTF_PT_0,
      O => FC1_CNT_2_RSTF
    );
  FC1_CNT_2_D1_528 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => FC1_CNT_2_D1
    );
  FC1_CNT_2_D2_PT_0_529 : X_AND2 
    port map (
      I0 => EXP14_EXP,
      I1 => EXP14_EXP,
      O => FC1_CNT_2_D2_PT_0
    );
  FC1_CNT_2_D2_PT_1_530 : X_AND4 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I1 => LIGHT_VALUE_5_FBK,
      I2 => LIGHT_VALUE_2_FBK,
      I3 => LIGHT_VALUE_3_FBK,
      O => FC1_CNT_2_D2_PT_1
    );
  FC1_CNT_2_D2_PT_2_531 : X_AND16 
    port map (
      I0 => FC1_CNT_2_D2_PT_2_0_INV,
      I1 => FC1_CNT_2_D2_PT_2_1_INV,
      I2 => FC1_CNT_2_D2_PT_2_2_INV,
      I3 => FC1_CNT_2_D2_PT_2_3_INV,
      I4 => FC1_CNT_2_D2_PT_2_4_INV,
      I5 => FC1_CNT_2_D2_PT_2_5_INV,
      I6 => FC1_CNT_2_D2_PT_2_6_INV,
      I7 => FC1_CNT_2_D2_PT_2_7_INV,
      I8 => FC1_CNT_2_D2_PT_2_8_INV,
      I9 => FC1_CNT_2_D2_PT_2_9_INV,
      I10 => FC1_CNT_2_D2_PT_2_10_INV,
      I11 => FC1_CNT_2_D2_PT_2_11_INV,
      I12 => FC1_CNT_2_D2_PT_2_12_INV,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_2_D2_PT_2
    );
  FC1_CNT_2_D2_532 : X_OR3 
    port map (
      I0 => FC1_CNT_2_D2_PT_0,
      I1 => FC1_CNT_2_D2_PT_1,
      I2 => FC1_CNT_2_D2_PT_2,
      O => FC1_CNT_2_D2
    );
  FC1_CNT_2_D_533 : X_XOR2 
    port map (
      I0 => FC1_CNT_2_D_TFF,
      I1 => FC1_CNT_2_Q,
      O => FC1_CNT_2_D
    );
  FC1_CNT_2_XOR : X_XOR2 
    port map (
      I0 => FC1_CNT_2_XOR_0_INV,
      I1 => FC1_CNT_2_D2,
      O => FC1_CNT_2_D_TFF
    );
  FC1_CNT_2_EXP_PT_0_534 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => FC1_CNT_2_EXP_PT_0_1_INV,
      I2 => FC1_CNT_2_EXP_PT_0_2_INV,
      I3 => FC1_CNT_2_EXP_PT_0_3_INV,
      I4 => FC1_CNT_2_EXP_PT_0_4_INV,
      I5 => FC1_CNT_2_EXP_PT_0_5_INV,
      I6 => FC1_CNT_2_EXP_PT_0_6_INV,
      I7 => FC1_CNT_2_EXP_PT_0_7_INV,
      I8 => FC1_CNT_2_EXP_PT_0_8_INV,
      I9 => FC1_CNT_2_EXP_PT_0_9_INV,
      I10 => LIGHT_VALUE_0_FBK,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_2_EXP_PT_0
    );
  FC1_CNT_2_EXP_PT_1_535 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => FC1_CNT_2_EXP_PT_1_1_INV,
      I2 => FC1_CNT_2_EXP_PT_1_2_INV,
      I3 => FC1_CNT_2_EXP_PT_1_3_INV,
      I4 => FC1_CNT_2_EXP_PT_1_4_INV,
      I5 => FC1_CNT_2_EXP_PT_1_5_INV,
      I6 => FC1_CNT_2_EXP_PT_1_6_INV,
      I7 => FC1_CNT_2_EXP_PT_1_7_INV,
      I8 => FC1_CNT_2_EXP_PT_1_8_INV,
      I9 => FC1_CNT_2_EXP_PT_1_9_INV,
      I10 => LIGHT_VALUE(4),
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_2_EXP_PT_1
    );
  FC1_CNT_2_EXP_536 : X_OR2 
    port map (
      I0 => FC1_CNT_2_EXP_PT_0,
      I1 => FC1_CNT_2_EXP_PT_1,
      O => FC1_CNT_2_EXP
    );
  FC1_CNT_2_FBK_537 : X_BUF 
    port map (
      I => FC1_CNT_2_Q,
      O => FC1_CNT_2_FBK
    );
  EXP14_EXP_PT_0_538 : X_AND2 
    port map (
      I0 => LIGHT_VALUE_1_EXP,
      I1 => LIGHT_VALUE_1_EXP,
      O => EXP14_EXP_PT_0
    );
  EXP14_EXP_PT_1_539 : X_AND2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => FC1_CNT_0_FBK,
      O => EXP14_EXP_PT_1
    );
  EXP14_EXP_PT_2_540 : X_AND2 
    port map (
      I0 => EXP14_EXP_PT_2_0_INV,
      I1 => EXP14_EXP_PT_2_1_INV,
      O => EXP14_EXP_PT_2
    );
  EXP14_EXP_PT_3_541 : X_AND2 
    port map (
      I0 => FC1_CNT_1_FBK,
      I1 => EXP14_EXP_PT_3_1_INV,
      O => EXP14_EXP_PT_3
    );
  EXP14_EXP_PT_4_542 : X_AND3 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I1 => LIGHT_VALUE_5_FBK,
      I2 => LIGHT_VALUE(4),
      O => EXP14_EXP_PT_4
    );
  EXP14_EXP_PT_5_543 : X_AND4 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I1 => LIGHT_VALUE_5_FBK,
      I2 => LIGHT_VALUE_1_FBK,
      I3 => LIGHT_VALUE_3_FBK,
      O => EXP14_EXP_PT_5
    );
  EXP14_EXP_544 : X_OR6 
    port map (
      I0 => EXP14_EXP_PT_0,
      I1 => EXP14_EXP_PT_1,
      I2 => EXP14_EXP_PT_2,
      I3 => EXP14_EXP_PT_3,
      I4 => EXP14_EXP_PT_4,
      I5 => EXP14_EXP_PT_5,
      O => EXP14_EXP
    );
  LIGHT_VALUE_1_Q_545 : X_BUF 
    port map (
      I => LIGHT_VALUE_1_Q,
      O => LIGHT_VALUE(1)
    );
  LIGHT_VALUE_1_REG : X_FF 
    port map (
      I => LIGHT_VALUE_1_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => LIGHT_VALUE_1_SETF,
      RST => PRLD,
      O => LIGHT_VALUE_1_Q
    );
  LIGHT_VALUE_1_SETF_PT_0_546 : X_AND2 
    port map (
      I0 => LIGHT_VALUE_1_SETF_PT_0_0_INV,
      I1 => LIGHT_VALUE_1_SETF_PT_0_1_INV,
      O => LIGHT_VALUE_1_SETF_PT_0
    );
  LIGHT_VALUE_1_SETF_547 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_1_SETF_PT_0,
      I1 => LIGHT_VALUE_1_SETF_PT_0,
      O => LIGHT_VALUE_1_SETF
    );
  LIGHT_VALUE_1_D1_548 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => LIGHT_VALUE_1_D1
    );
  LIGHT_VALUE_1_D2_PT_0_549 : X_AND2 
    port map (
      I0 => EXP13_EXP,
      I1 => EXP13_EXP,
      O => LIGHT_VALUE_1_D2_PT_0
    );
  LIGHT_VALUE_1_D2_PT_1_550 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => LIGHT_VALUE_1_D2_PT_1_1_INV,
      I2 => LIGHT_VALUE_1_D2_PT_1_2_INV,
      I3 => LIGHT_VALUE_1_D2_PT_1_3_INV,
      I4 => LIGHT_VALUE_1_D2_PT_1_4_INV,
      I5 => LIGHT_VALUE_1_D2_PT_1_5_INV,
      I6 => LIGHT_VALUE_1_D2_PT_1_6_INV,
      I7 => LIGHT_VALUE_1_D2_PT_1_7_INV,
      I8 => LIGHT_VALUE_1_D2_PT_1_8_INV,
      I9 => LIGHT_VALUE_1_D2_PT_1_9_INV,
      I10 => LIGHT_VALUE_1_FBK,
      I11 => LIGHT_VALUE_1_D2_PT_1_11_INV,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_1_D2_PT_1
    );
  LIGHT_VALUE_1_D2_PT_2_551 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => LIGHT_VALUE_1_D2_PT_2_1_INV,
      I2 => LIGHT_VALUE_1_D2_PT_2_2_INV,
      I3 => LIGHT_VALUE_1_D2_PT_2_3_INV,
      I4 => LIGHT_VALUE_1_D2_PT_2_4_INV,
      I5 => LIGHT_VALUE_1_D2_PT_2_5_INV,
      I6 => LIGHT_VALUE_1_D2_PT_2_6_INV,
      I7 => LIGHT_VALUE_1_D2_PT_2_7_INV,
      I8 => LIGHT_VALUE_1_D2_PT_2_8_INV,
      I9 => LIGHT_VALUE_1_D2_PT_2_9_INV,
      I10 => LIGHT_VALUE_2_FBK,
      I11 => LIGHT_VALUE_1_D2_PT_2_11_INV,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_1_D2_PT_2
    );
  LIGHT_VALUE_1_D2_PT_3_552 : X_AND16 
    port map (
      I0 => LIGHT_VALUE_1_D2_PT_3_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I2 => LIGHT_VALUE_1_D2_PT_3_2_INV,
      I3 => FC1_CNT_1_FBK,
      I4 => FC1_CNT_2_FBK,
      I5 => FC1_CNT_0_FBK,
      I6 => FC1_CNT(3),
      I7 => FC1_CNT(4),
      I8 => FC1_CNT(5),
      I9 => FC1_CNT(6),
      I10 => FC1_CNT(7),
      I11 => LIGHT_VALUE_0_FBK,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_1_D2_PT_3
    );
  LIGHT_VALUE_1_D2_553 : X_OR4 
    port map (
      I0 => LIGHT_VALUE_1_D2_PT_0,
      I1 => LIGHT_VALUE_1_D2_PT_1,
      I2 => LIGHT_VALUE_1_D2_PT_2,
      I3 => LIGHT_VALUE_1_D2_PT_3,
      O => LIGHT_VALUE_1_D2
    );
  LIGHT_VALUE_1_D_554 : X_XOR2 
    port map (
      I0 => LIGHT_VALUE_1_D_TFF,
      I1 => LIGHT_VALUE_1_Q,
      O => LIGHT_VALUE_1_D
    );
  LIGHT_VALUE_1_XOR : X_XOR2 
    port map (
      I0 => LIGHT_VALUE_1_D1,
      I1 => LIGHT_VALUE_1_D2,
      O => LIGHT_VALUE_1_D_TFF
    );
  LIGHT_VALUE_1_EXP_PT_0_555 : X_AND2 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I1 => LIGHT_VALUE_1_EXP_PT_0_1_INV,
      O => LIGHT_VALUE_1_EXP_PT_0
    );
  LIGHT_VALUE_1_EXP_556 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_1_EXP_PT_0,
      I1 => LIGHT_VALUE_1_EXP_PT_0,
      O => LIGHT_VALUE_1_EXP
    );
  LIGHT_VALUE_1_FBK_557 : X_BUF 
    port map (
      I => LIGHT_VALUE_1_Q,
      O => LIGHT_VALUE_1_FBK
    );
  EXP13_EXP_PT_0_558 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => EXP13_EXP_PT_0_1_INV,
      I2 => LIGHT_VALUE_5_FBK,
      I3 => EXP13_EXP_PT_0_3_INV,
      I4 => EXP13_EXP_PT_0_4_INV,
      I5 => EXP13_EXP_PT_0_5_INV,
      I6 => EXP13_EXP_PT_0_6_INV,
      I7 => EXP13_EXP_PT_0_7_INV,
      I8 => EXP13_EXP_PT_0_8_INV,
      I9 => EXP13_EXP_PT_0_9_INV,
      I10 => EXP13_EXP_PT_0_10_INV,
      I11 => EXP13_EXP_PT_0_11_INV,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP13_EXP_PT_0
    );
  EXP13_EXP_PT_1_559 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => EXP13_EXP_PT_1_1_INV,
      I2 => EXP13_EXP_PT_1_2_INV,
      I3 => EXP13_EXP_PT_1_3_INV,
      I4 => EXP13_EXP_PT_1_4_INV,
      I5 => EXP13_EXP_PT_1_5_INV,
      I6 => EXP13_EXP_PT_1_6_INV,
      I7 => EXP13_EXP_PT_1_7_INV,
      I8 => EXP13_EXP_PT_1_8_INV,
      I9 => EXP13_EXP_PT_1_9_INV,
      I10 => EXP13_EXP_PT_1_10_INV,
      I11 => LIGHT_VALUE_3_FBK,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP13_EXP_PT_1
    );
  EXP13_EXP_PT_2_560 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => EXP13_EXP_PT_2_1_INV,
      I2 => EXP13_EXP_PT_2_2_INV,
      I3 => EXP13_EXP_PT_2_3_INV,
      I4 => EXP13_EXP_PT_2_4_INV,
      I5 => EXP13_EXP_PT_2_5_INV,
      I6 => EXP13_EXP_PT_2_6_INV,
      I7 => EXP13_EXP_PT_2_7_INV,
      I8 => EXP13_EXP_PT_2_8_INV,
      I9 => EXP13_EXP_PT_2_9_INV,
      I10 => EXP13_EXP_PT_2_10_INV,
      I11 => LIGHT_VALUE(4),
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP13_EXP_PT_2
    );
  EXP13_EXP_PT_3_561 : X_AND16 
    port map (
      I0 => EXP13_EXP_PT_3_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I2 => FC1_CNT_1_FBK,
      I3 => FC1_CNT_2_FBK,
      I4 => FC1_CNT_0_FBK,
      I5 => FC1_CNT(3),
      I6 => FC1_CNT(4),
      I7 => FC1_CNT(5),
      I8 => FC1_CNT(6),
      I9 => FC1_CNT(7),
      I10 => LIGHT_VALUE_0_FBK,
      I11 => EXP13_EXP_PT_3_11_INV,
      I12 => EXP13_EXP_PT_3_12_INV,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP13_EXP_PT_3
    );
  EXP13_EXP_PT_4_562 : X_AND16 
    port map (
      I0 => EXP13_EXP_PT_4_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I2 => FC1_CNT_1_FBK,
      I3 => FC1_CNT_2_FBK,
      I4 => FC1_CNT_0_FBK,
      I5 => FC1_CNT(3),
      I6 => FC1_CNT(4),
      I7 => FC1_CNT(5),
      I8 => FC1_CNT(6),
      I9 => FC1_CNT(7),
      I10 => EXP13_EXP_PT_4_10_INV,
      I11 => EXP13_EXP_PT_4_11_INV,
      I12 => LIGHT_VALUE_0_FBK,
      I13 => EXP13_EXP_PT_4_13_INV,
      I14 => VCC,
      I15 => VCC,
      O => EXP13_EXP_PT_4
    );
  EXP13_EXP_563 : X_OR5 
    port map (
      I0 => EXP13_EXP_PT_0,
      I1 => EXP13_EXP_PT_1,
      I2 => EXP13_EXP_PT_2,
      I3 => EXP13_EXP_PT_3,
      I4 => EXP13_EXP_PT_4,
      O => EXP13_EXP
    );
  FC1_CNT_4_Q_564 : X_BUF 
    port map (
      I => FC1_CNT_4_Q,
      O => FC1_CNT(4)
    );
  FC1_CNT_4_R_OR_PRLD_565 : X_OR2 
    port map (
      I0 => FC1_CNT_4_RSTF,
      I1 => PRLD,
      O => FC1_CNT_4_R_OR_PRLD
    );
  FC1_CNT_4_REG : X_FF 
    port map (
      I => FC1_CNT_4_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => FC1_CNT_4_R_OR_PRLD,
      O => FC1_CNT_4_Q
    );
  FC1_CNT_4_RSTF_PT_0_566 : X_AND2 
    port map (
      I0 => FC1_CNT_4_RSTF_PT_0_0_INV,
      I1 => FC1_CNT_4_RSTF_PT_0_1_INV,
      O => FC1_CNT_4_RSTF_PT_0
    );
  FC1_CNT_4_RSTF_567 : X_OR2 
    port map (
      I0 => FC1_CNT_4_RSTF_PT_0,
      I1 => FC1_CNT_4_RSTF_PT_0,
      O => FC1_CNT_4_RSTF
    );
  FC1_CNT_4_D1_568 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => FC1_CNT_4_D1
    );
  FC1_CNT_4_D2_PT_0_569 : X_AND2 
    port map (
      I0 => LIGHT_VALUE_4_EXP,
      I1 => LIGHT_VALUE_4_EXP,
      O => FC1_CNT_4_D2_PT_0
    );
  FC1_CNT_4_D2_PT_1_570 : X_AND2 
    port map (
      I0 => EXP8_EXP,
      I1 => EXP8_EXP,
      O => FC1_CNT_4_D2_PT_1
    );
  FC1_CNT_4_D2_PT_2_571 : X_AND7 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => FC1_CNT_3_FBK,
      I2 => FC1_CNT(1),
      I3 => FC1_CNT(2),
      I4 => FC1_CNT(0),
      I5 => FC1_CNT_4_D2_PT_2_5_INV,
      I6 => FC1_CNT_4_D2_PT_2_6_INV,
      O => FC1_CNT_4_D2_PT_2
    );
  FC1_CNT_4_D2_PT_3_572 : X_AND7 
    port map (
      I0 => FC1_CNT_4_D2_PT_3_0_INV,
      I1 => FC1_CNT_4_D2_PT_3_1_INV,
      I2 => FC1_CNT_4_D2_PT_3_2_INV,
      I3 => FC1_CNT_4_D2_PT_3_3_INV,
      I4 => FC1_CNT_4_FBK,
      I5 => FC1_CNT_4_D2_PT_3_5_INV,
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_4_D2_PT_3
    );
  FC1_CNT_4_D2_PT_4_573 : X_AND7 
    port map (
      I0 => FC1_CNT_4_D2_PT_4_0_INV,
      I1 => FC1_CNT_4_D2_PT_4_1_INV,
      I2 => FC1_CNT_4_D2_PT_4_2_INV,
      I3 => FC1_CNT_4_D2_PT_4_3_INV,
      I4 => FC1_CNT_6_FBK,
      I5 => FC1_CNT_4_D2_PT_4_5_INV,
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_4_D2_PT_4
    );
  FC1_CNT_4_D2_PT_5_574 : X_AND7 
    port map (
      I0 => FC1_CNT_4_D2_PT_5_0_INV,
      I1 => FC1_CNT_4_D2_PT_5_1_INV,
      I2 => FC1_CNT_4_D2_PT_5_2_INV,
      I3 => FC1_CNT_4_D2_PT_5_3_INV,
      I4 => FC1_CNT_4_D2_PT_5_4_INV,
      I5 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I6 => FC1_CNT_7_FBK,
      O => FC1_CNT_4_D2_PT_5
    );
  FC1_CNT_4_D2_575 : X_OR6 
    port map (
      I0 => FC1_CNT_4_D2_PT_0,
      I1 => FC1_CNT_4_D2_PT_1,
      I2 => FC1_CNT_4_D2_PT_2,
      I3 => FC1_CNT_4_D2_PT_3,
      I4 => FC1_CNT_4_D2_PT_4,
      I5 => FC1_CNT_4_D2_PT_5,
      O => FC1_CNT_4_D2
    );
  FC1_CNT_4_D_576 : X_XOR2 
    port map (
      I0 => FC1_CNT_4_D_TFF,
      I1 => FC1_CNT_4_Q,
      O => FC1_CNT_4_D
    );
  FC1_CNT_4_XOR : X_XOR2 
    port map (
      I0 => FC1_CNT_4_D1,
      I1 => FC1_CNT_4_D2,
      O => FC1_CNT_4_D_TFF
    );
  FC1_CNT_4_FBK_577 : X_BUF 
    port map (
      I => FC1_CNT_4_Q,
      O => FC1_CNT_4_FBK
    );
  EXP8_EXP_PT_0_578 : X_AND2 
    port map (
      I0 => FC1_CNT_5_EXP,
      I1 => FC1_CNT_5_EXP,
      O => EXP8_EXP_PT_0
    );
  EXP8_EXP_PT_1_579 : X_AND7 
    port map (
      I0 => EXP8_EXP_PT_1_0_INV,
      I1 => EXP8_EXP_PT_1_1_INV,
      I2 => EXP8_EXP_PT_1_2_INV,
      I3 => EXP8_EXP_PT_1_3_INV,
      I4 => FC1_CNT_5_FBK,
      I5 => EXP8_EXP_PT_1_5_INV,
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP8_EXP_PT_1
    );
  EXP8_EXP_PT_2_580 : X_AND7 
    port map (
      I0 => EXP8_EXP_PT_2_0_INV,
      I1 => EXP8_EXP_PT_2_1_INV,
      I2 => EXP8_EXP_PT_2_2_INV,
      I3 => EXP8_EXP_PT_2_3_INV,
      I4 => EXP8_EXP_PT_2_4_INV,
      I5 => LIGHT_VALUE(3),
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP8_EXP_PT_2
    );
  EXP8_EXP_PT_3_581 : X_AND7 
    port map (
      I0 => EXP8_EXP_PT_3_0_INV,
      I1 => EXP8_EXP_PT_3_1_INV,
      I2 => EXP8_EXP_PT_3_2_INV,
      I3 => EXP8_EXP_PT_3_3_INV,
      I4 => EXP8_EXP_PT_3_4_INV,
      I5 => LIGHT_VALUE(1),
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP8_EXP_PT_3
    );
  EXP8_EXP_PT_4_582 : X_AND7 
    port map (
      I0 => EXP8_EXP_PT_4_0_INV,
      I1 => EXP8_EXP_PT_4_1_INV,
      I2 => EXP8_EXP_PT_4_2_INV,
      I3 => EXP8_EXP_PT_4_3_INV,
      I4 => EXP8_EXP_PT_4_4_INV,
      I5 => LIGHT_VALUE(2),
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP8_EXP_PT_4
    );
  EXP8_EXP_PT_5_583 : X_AND7 
    port map (
      I0 => EXP8_EXP_PT_5_0_INV,
      I1 => EXP8_EXP_PT_5_1_INV,
      I2 => EXP8_EXP_PT_5_2_INV,
      I3 => EXP8_EXP_PT_5_3_INV,
      I4 => EXP8_EXP_PT_5_4_INV,
      I5 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I6 => LIGHT_VALUE(0),
      O => EXP8_EXP_PT_5
    );
  EXP8_EXP_584 : X_OR6 
    port map (
      I0 => EXP8_EXP_PT_0,
      I1 => EXP8_EXP_PT_1,
      I2 => EXP8_EXP_PT_2,
      I3 => EXP8_EXP_PT_3,
      I4 => EXP8_EXP_PT_4,
      I5 => EXP8_EXP_PT_5,
      O => EXP8_EXP
    );
  FC1_CNT_5_Q_585 : X_BUF 
    port map (
      I => FC1_CNT_5_Q,
      O => FC1_CNT(5)
    );
  FC1_CNT_5_R_OR_PRLD_586 : X_OR2 
    port map (
      I0 => FC1_CNT_5_RSTF,
      I1 => PRLD,
      O => FC1_CNT_5_R_OR_PRLD
    );
  FC1_CNT_5_REG : X_FF 
    port map (
      I => FC1_CNT_5_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => FC1_CNT_5_R_OR_PRLD,
      O => FC1_CNT_5_Q
    );
  FC1_CNT_5_RSTF_PT_0_587 : X_AND2 
    port map (
      I0 => FC1_CNT_5_RSTF_PT_0_0_INV,
      I1 => FC1_CNT_5_RSTF_PT_0_1_INV,
      O => FC1_CNT_5_RSTF_PT_0
    );
  FC1_CNT_5_RSTF_588 : X_OR2 
    port map (
      I0 => FC1_CNT_5_RSTF_PT_0,
      I1 => FC1_CNT_5_RSTF_PT_0,
      O => FC1_CNT_5_RSTF
    );
  FC1_CNT_5_D1_589 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => FC1_CNT_5_D1
    );
  FC1_CNT_5_D2_PT_0_590 : X_AND2 
    port map (
      I0 => EXP7_EXP,
      I1 => EXP7_EXP,
      O => FC1_CNT_5_D2_PT_0
    );
  FC1_CNT_5_D2_PT_1_591 : X_AND8 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => FC1_CNT_3_FBK,
      I2 => FC1_CNT(1),
      I3 => FC1_CNT(2),
      I4 => FC1_CNT_4_FBK,
      I5 => FC1_CNT(0),
      I6 => FC1_CNT_5_D2_PT_1_6_INV,
      I7 => FC1_CNT_5_D2_PT_1_7_INV,
      O => FC1_CNT_5_D2_PT_1
    );
  FC1_CNT_5_D2_PT_2_592 : X_AND8 
    port map (
      I0 => FC1_CNT_5_D2_PT_2_0_INV,
      I1 => FC1_CNT_5_D2_PT_2_1_INV,
      I2 => FC1_CNT_5_D2_PT_2_2_INV,
      I3 => FC1_CNT_5_D2_PT_2_3_INV,
      I4 => FC1_CNT_5_D2_PT_2_4_INV,
      I5 => FC1_CNT_6_FBK,
      I6 => FC1_CNT_5_D2_PT_2_6_INV,
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_5_D2_PT_2
    );
  FC1_CNT_5_D2_PT_3_593 : X_AND8 
    port map (
      I0 => FC1_CNT_5_D2_PT_3_0_INV,
      I1 => FC1_CNT_5_D2_PT_3_1_INV,
      I2 => FC1_CNT_5_D2_PT_3_2_INV,
      I3 => FC1_CNT_5_D2_PT_3_3_INV,
      I4 => FC1_CNT_5_D2_PT_3_4_INV,
      I5 => FC1_CNT_5_D2_PT_3_5_INV,
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I7 => FC1_CNT_7_FBK,
      O => FC1_CNT_5_D2_PT_3
    );
  FC1_CNT_5_D2_594 : X_OR4 
    port map (
      I0 => FC1_CNT_5_D2_PT_0,
      I1 => FC1_CNT_5_D2_PT_1,
      I2 => FC1_CNT_5_D2_PT_2,
      I3 => FC1_CNT_5_D2_PT_3,
      O => FC1_CNT_5_D2
    );
  FC1_CNT_5_D_595 : X_XOR2 
    port map (
      I0 => FC1_CNT_5_D_TFF,
      I1 => FC1_CNT_5_Q,
      O => FC1_CNT_5_D
    );
  FC1_CNT_5_XOR : X_XOR2 
    port map (
      I0 => FC1_CNT_5_D1,
      I1 => FC1_CNT_5_D2,
      O => FC1_CNT_5_D_TFF
    );
  FC1_CNT_5_EXP_PT_0_596 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => FC1_CNT_5_EXP_PT_0_1_INV,
      I2 => FC1_CNT_3_FBK,
      I3 => FC1_CNT(1),
      I4 => FC1_CNT(2),
      I5 => FC1_CNT(0),
      I6 => FC1_CNT_5_EXP_PT_0_6_INV,
      I7 => FC1_CNT_5_EXP_PT_0_7_INV,
      I8 => FC1_CNT_5_EXP_PT_0_8_INV,
      I9 => VCC,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_5_EXP_PT_0
    );
  FC1_CNT_5_EXP_597 : X_OR2 
    port map (
      I0 => FC1_CNT_5_EXP_PT_0,
      I1 => FC1_CNT_5_EXP_PT_0,
      O => FC1_CNT_5_EXP
    );
  FC1_CNT_5_FBK_598 : X_BUF 
    port map (
      I => FC1_CNT_5_Q,
      O => FC1_CNT_5_FBK
    );
  EXP7_EXP_PT_0_599 : X_AND2 
    port map (
      I0 => EXP6_EXP,
      I1 => EXP6_EXP,
      O => EXP7_EXP_PT_0
    );
  EXP7_EXP_PT_1_600 : X_AND8 
    port map (
      I0 => EXP7_EXP_PT_1_0_INV,
      I1 => EXP7_EXP_PT_1_1_INV,
      I2 => EXP7_EXP_PT_1_2_INV,
      I3 => EXP7_EXP_PT_1_3_INV,
      I4 => EXP7_EXP_PT_1_4_INV,
      I5 => FC1_CNT_5_FBK,
      I6 => EXP7_EXP_PT_1_6_INV,
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP7_EXP_PT_1
    );
  EXP7_EXP_PT_2_601 : X_AND8 
    port map (
      I0 => EXP7_EXP_PT_2_0_INV,
      I1 => EXP7_EXP_PT_2_1_INV,
      I2 => EXP7_EXP_PT_2_2_INV,
      I3 => EXP7_EXP_PT_2_3_INV,
      I4 => EXP7_EXP_PT_2_4_INV,
      I5 => EXP7_EXP_PT_2_5_INV,
      I6 => LIGHT_VALUE(3),
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP7_EXP_PT_2
    );
  EXP7_EXP_PT_3_602 : X_AND8 
    port map (
      I0 => EXP7_EXP_PT_3_0_INV,
      I1 => EXP7_EXP_PT_3_1_INV,
      I2 => EXP7_EXP_PT_3_2_INV,
      I3 => EXP7_EXP_PT_3_3_INV,
      I4 => EXP7_EXP_PT_3_4_INV,
      I5 => EXP7_EXP_PT_3_5_INV,
      I6 => LIGHT_VALUE(1),
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP7_EXP_PT_3
    );
  EXP7_EXP_PT_4_603 : X_AND8 
    port map (
      I0 => EXP7_EXP_PT_4_0_INV,
      I1 => EXP7_EXP_PT_4_1_INV,
      I2 => EXP7_EXP_PT_4_2_INV,
      I3 => EXP7_EXP_PT_4_3_INV,
      I4 => EXP7_EXP_PT_4_4_INV,
      I5 => EXP7_EXP_PT_4_5_INV,
      I6 => LIGHT_VALUE(2),
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP7_EXP_PT_4
    );
  EXP7_EXP_PT_5_604 : X_AND8 
    port map (
      I0 => EXP7_EXP_PT_5_0_INV,
      I1 => EXP7_EXP_PT_5_1_INV,
      I2 => EXP7_EXP_PT_5_2_INV,
      I3 => EXP7_EXP_PT_5_3_INV,
      I4 => EXP7_EXP_PT_5_4_INV,
      I5 => EXP7_EXP_PT_5_5_INV,
      I6 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I7 => LIGHT_VALUE(0),
      O => EXP7_EXP_PT_5
    );
  EXP7_EXP_605 : X_OR6 
    port map (
      I0 => EXP7_EXP_PT_0,
      I1 => EXP7_EXP_PT_1,
      I2 => EXP7_EXP_PT_2,
      I3 => EXP7_EXP_PT_3,
      I4 => EXP7_EXP_PT_4,
      I5 => EXP7_EXP_PT_5,
      O => EXP7_EXP
    );
  EXP6_EXP_PT_0_606 : X_AND8 
    port map (
      I0 => EXP6_EXP_PT_0_0_INV,
      I1 => LIGHT_VALUE_4_FBK,
      I2 => EXP6_EXP_PT_0_2_INV,
      I3 => EXP6_EXP_PT_0_3_INV,
      I4 => EXP6_EXP_PT_0_4_INV,
      I5 => EXP6_EXP_PT_0_5_INV,
      I6 => EXP6_EXP_PT_0_6_INV,
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP6_EXP_PT_0
    );
  EXP6_EXP_PT_1_607 : X_AND8 
    port map (
      I0 => EXP6_EXP_PT_1_0_INV,
      I1 => EXP6_EXP_PT_1_1_INV,
      I2 => EXP6_EXP_PT_1_2_INV,
      I3 => EXP6_EXP_PT_1_3_INV,
      I4 => EXP6_EXP_PT_1_4_INV,
      I5 => EXP6_EXP_PT_1_5_INV,
      I6 => LIGHT_VALUE(5),
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP6_EXP_PT_1
    );
  EXP6_EXP_PT_2_608 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => EXP6_EXP_PT_2_1_INV,
      I2 => FC1_CNT_3_FBK,
      I3 => FC1_CNT(1),
      I4 => FC1_CNT(2),
      I5 => FC1_CNT_4_FBK,
      I6 => FC1_CNT(0),
      I7 => EXP6_EXP_PT_2_7_INV,
      I8 => EXP6_EXP_PT_2_8_INV,
      I9 => VCC,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP6_EXP_PT_2
    );
  EXP6_EXP_PT_3_609 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => EXP6_EXP_PT_3_1_INV,
      I2 => FC1_CNT_3_FBK,
      I3 => FC1_CNT(1),
      I4 => FC1_CNT(2),
      I5 => FC1_CNT_4_FBK,
      I6 => FC1_CNT(0),
      I7 => EXP6_EXP_PT_3_7_INV,
      I8 => EXP6_EXP_PT_3_8_INV,
      I9 => EXP6_EXP_PT_3_9_INV,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP6_EXP_PT_3
    );
  EXP6_EXP_610 : X_OR4 
    port map (
      I0 => EXP6_EXP_PT_0,
      I1 => EXP6_EXP_PT_1,
      I2 => EXP6_EXP_PT_2,
      I3 => EXP6_EXP_PT_3,
      O => EXP6_EXP
    );
  LIGHT_VALUE_3_Q_611 : X_BUF 
    port map (
      I => LIGHT_VALUE_3_Q,
      O => LIGHT_VALUE(3)
    );
  LIGHT_VALUE_3_REG : X_FF 
    port map (
      I => LIGHT_VALUE_3_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => LIGHT_VALUE_3_SETF,
      RST => PRLD,
      O => LIGHT_VALUE_3_Q
    );
  LIGHT_VALUE_3_SETF_PT_0_612 : X_AND2 
    port map (
      I0 => LIGHT_VALUE_3_SETF_PT_0_0_INV,
      I1 => LIGHT_VALUE_3_SETF_PT_0_1_INV,
      O => LIGHT_VALUE_3_SETF_PT_0
    );
  LIGHT_VALUE_3_SETF_613 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_3_SETF_PT_0,
      I1 => LIGHT_VALUE_3_SETF_PT_0,
      O => LIGHT_VALUE_3_SETF
    );
  LIGHT_VALUE_3_D1_614 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => LIGHT_VALUE_3_D1
    );
  LIGHT_VALUE_3_D2_PT_0_615 : X_AND2 
    port map (
      I0 => LIGHT_VALUE_5_EXP,
      I1 => LIGHT_VALUE_5_EXP,
      O => LIGHT_VALUE_3_D2_PT_0
    );
  LIGHT_VALUE_3_D2_PT_1_616 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => LIGHT_VALUE_3_D2_PT_1_1_INV,
      I2 => LIGHT_VALUE_3_D2_PT_1_2_INV,
      I3 => LIGHT_VALUE_3_D2_PT_1_3_INV,
      I4 => LIGHT_VALUE_3_D2_PT_1_4_INV,
      I5 => LIGHT_VALUE_3_D2_PT_1_5_INV,
      I6 => LIGHT_VALUE_3_D2_PT_1_6_INV,
      I7 => LIGHT_VALUE_3_D2_PT_1_7_INV,
      I8 => LIGHT_VALUE_3_D2_PT_1_8_INV,
      I9 => LIGHT_VALUE_3_D2_PT_1_9_INV,
      I10 => LIGHT_VALUE_3_D2_PT_1_10_INV,
      I11 => LIGHT_VALUE_3_D2_PT_1_11_INV,
      I12 => LIGHT_VALUE_3_D2_PT_1_12_INV,
      I13 => LIGHT_VALUE_3_FBK,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_3_D2_PT_1
    );
  LIGHT_VALUE_3_D2_PT_2_617 : X_AND16 
    port map (
      I0 => LIGHT_VALUE_3_D2_PT_2_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I2 => LIGHT_VALUE_3_D2_PT_2_2_INV,
      I3 => FC1_CNT_1_FBK,
      I4 => FC1_CNT_2_FBK,
      I5 => FC1_CNT_0_FBK,
      I6 => FC1_CNT(3),
      I7 => FC1_CNT(4),
      I8 => FC1_CNT(5),
      I9 => FC1_CNT(6),
      I10 => FC1_CNT(7),
      I11 => LIGHT_VALUE_1_FBK,
      I12 => LIGHT_VALUE_2_FBK,
      I13 => LIGHT_VALUE_0_FBK,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_3_D2_PT_2
    );
  LIGHT_VALUE_3_D2_618 : X_OR3 
    port map (
      I0 => LIGHT_VALUE_3_D2_PT_0,
      I1 => LIGHT_VALUE_3_D2_PT_1,
      I2 => LIGHT_VALUE_3_D2_PT_2,
      O => LIGHT_VALUE_3_D2
    );
  LIGHT_VALUE_3_D_619 : X_XOR2 
    port map (
      I0 => LIGHT_VALUE_3_D_TFF,
      I1 => LIGHT_VALUE_3_Q,
      O => LIGHT_VALUE_3_D
    );
  LIGHT_VALUE_3_XOR : X_XOR2 
    port map (
      I0 => LIGHT_VALUE_3_D1,
      I1 => LIGHT_VALUE_3_D2,
      O => LIGHT_VALUE_3_D_TFF
    );
  LIGHT_VALUE_3_EXP_PT_0_620 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => LIGHT_VALUE_3_EXP_PT_0_1_INV,
      I2 => LIGHT_VALUE_5_FBK,
      I3 => LIGHT_VALUE_3_EXP_PT_0_3_INV,
      I4 => LIGHT_VALUE_3_EXP_PT_0_4_INV,
      I5 => LIGHT_VALUE_3_EXP_PT_0_5_INV,
      I6 => LIGHT_VALUE_3_EXP_PT_0_6_INV,
      I7 => LIGHT_VALUE_3_EXP_PT_0_7_INV,
      I8 => LIGHT_VALUE_3_EXP_PT_0_8_INV,
      I9 => LIGHT_VALUE_3_EXP_PT_0_9_INV,
      I10 => LIGHT_VALUE_3_EXP_PT_0_10_INV,
      I11 => LIGHT_VALUE_3_EXP_PT_0_11_INV,
      I12 => LIGHT_VALUE_3_EXP_PT_0_12_INV,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_3_EXP_PT_0
    );
  LIGHT_VALUE_3_EXP_PT_1_621 : X_AND16 
    port map (
      I0 => LIGHT_VALUE_3_EXP_PT_1_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I2 => FC1_CNT_1_FBK,
      I3 => FC1_CNT_2_FBK,
      I4 => FC1_CNT_0_FBK,
      I5 => FC1_CNT(3),
      I6 => FC1_CNT(4),
      I7 => FC1_CNT(5),
      I8 => FC1_CNT(6),
      I9 => FC1_CNT(7),
      I10 => LIGHT_VALUE_1_FBK,
      I11 => LIGHT_VALUE_0_FBK,
      I12 => LIGHT_VALUE_3_EXP_PT_1_12_INV,
      I13 => LIGHT_VALUE_3_EXP_PT_1_13_INV,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_3_EXP_PT_1
    );
  LIGHT_VALUE_3_EXP_622 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_3_EXP_PT_0,
      I1 => LIGHT_VALUE_3_EXP_PT_1,
      O => LIGHT_VALUE_3_EXP
    );
  LIGHT_VALUE_3_FBK_623 : X_BUF 
    port map (
      I => LIGHT_VALUE_3_Q,
      O => LIGHT_VALUE_3_FBK
    );
  FC1_CNT_6_Q_624 : X_BUF 
    port map (
      I => FC1_CNT_6_Q,
      O => FC1_CNT(6)
    );
  FC1_CNT_6_R_OR_PRLD_625 : X_OR2 
    port map (
      I0 => FC1_CNT_6_RSTF,
      I1 => PRLD,
      O => FC1_CNT_6_R_OR_PRLD
    );
  FC1_CNT_6_REG : X_FF 
    port map (
      I => FC1_CNT_6_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => FC1_CNT_6_R_OR_PRLD,
      O => FC1_CNT_6_Q
    );
  FC1_CNT_6_RSTF_PT_0_626 : X_AND2 
    port map (
      I0 => FC1_CNT_6_RSTF_PT_0_0_INV,
      I1 => FC1_CNT_6_RSTF_PT_0_1_INV,
      O => FC1_CNT_6_RSTF_PT_0
    );
  FC1_CNT_6_RSTF_627 : X_OR2 
    port map (
      I0 => FC1_CNT_6_RSTF_PT_0,
      I1 => FC1_CNT_6_RSTF_PT_0,
      O => FC1_CNT_6_RSTF
    );
  FC1_CNT_6_D1_628 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => FC1_CNT_6_D1
    );
  FC1_CNT_6_D2_PT_0_629 : X_AND2 
    port map (
      I0 => FC1_CNT_3_EXP,
      I1 => FC1_CNT_3_EXP,
      O => FC1_CNT_6_D2_PT_0
    );
  FC1_CNT_6_D2_PT_1_630 : X_AND2 
    port map (
      I0 => EXP5_EXP,
      I1 => EXP5_EXP,
      O => FC1_CNT_6_D2_PT_1
    );
  FC1_CNT_6_D2_PT_2_631 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => FC1_CNT_3_FBK,
      I2 => FC1_CNT(1),
      I3 => FC1_CNT(2),
      I4 => FC1_CNT_4_FBK,
      I5 => FC1_CNT_5_FBK,
      I6 => FC1_CNT(0),
      I7 => FC1_CNT_6_D2_PT_2_7_INV,
      I8 => FC1_CNT_6_D2_PT_2_8_INV,
      I9 => VCC,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_6_D2_PT_2
    );
  FC1_CNT_6_D2_PT_3_632 : X_AND16 
    port map (
      I0 => FC1_CNT_6_D2_PT_3_0_INV,
      I1 => FC1_CNT_6_D2_PT_3_1_INV,
      I2 => FC1_CNT_6_D2_PT_3_2_INV,
      I3 => FC1_CNT_6_D2_PT_3_3_INV,
      I4 => FC1_CNT_6_D2_PT_3_4_INV,
      I5 => FC1_CNT_6_D2_PT_3_5_INV,
      I6 => FC1_CNT_6_FBK,
      I7 => FC1_CNT_6_D2_PT_3_7_INV,
      I8 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I9 => VCC,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_6_D2_PT_3
    );
  FC1_CNT_6_D2_PT_4_633 : X_AND16 
    port map (
      I0 => FC1_CNT_6_D2_PT_4_0_INV,
      I1 => FC1_CNT_6_D2_PT_4_1_INV,
      I2 => FC1_CNT_6_D2_PT_4_2_INV,
      I3 => FC1_CNT_6_D2_PT_4_3_INV,
      I4 => FC1_CNT_6_D2_PT_4_4_INV,
      I5 => FC1_CNT_6_D2_PT_4_5_INV,
      I6 => FC1_CNT_6_D2_PT_4_6_INV,
      I7 => LIGHT_VALUE(2),
      I8 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I9 => VCC,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_6_D2_PT_4
    );
  FC1_CNT_6_D2_PT_5_634 : X_AND16 
    port map (
      I0 => FC1_CNT_6_D2_PT_5_0_INV,
      I1 => FC1_CNT_6_D2_PT_5_1_INV,
      I2 => FC1_CNT_6_D2_PT_5_2_INV,
      I3 => FC1_CNT_6_D2_PT_5_3_INV,
      I4 => FC1_CNT_6_D2_PT_5_4_INV,
      I5 => FC1_CNT_6_D2_PT_5_5_INV,
      I6 => FC1_CNT_6_D2_PT_5_6_INV,
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I8 => FC1_CNT_7_FBK,
      I9 => VCC,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => FC1_CNT_6_D2_PT_5
    );
  FC1_CNT_6_D2_635 : X_OR6 
    port map (
      I0 => FC1_CNT_6_D2_PT_0,
      I1 => FC1_CNT_6_D2_PT_1,
      I2 => FC1_CNT_6_D2_PT_2,
      I3 => FC1_CNT_6_D2_PT_3,
      I4 => FC1_CNT_6_D2_PT_4,
      I5 => FC1_CNT_6_D2_PT_5,
      O => FC1_CNT_6_D2
    );
  FC1_CNT_6_D_636 : X_XOR2 
    port map (
      I0 => FC1_CNT_6_D_TFF,
      I1 => FC1_CNT_6_Q,
      O => FC1_CNT_6_D
    );
  FC1_CNT_6_XOR : X_XOR2 
    port map (
      I0 => FC1_CNT_6_D1,
      I1 => FC1_CNT_6_D2,
      O => FC1_CNT_6_D_TFF
    );
  FC1_CNT_6_FBK_637 : X_BUF 
    port map (
      I => FC1_CNT_6_Q,
      O => FC1_CNT_6_FBK
    );
  EXP5_EXP_PT_0_638 : X_AND16 
    port map (
      I0 => EXP5_EXP_PT_0_0_INV,
      I1 => LIGHT_VALUE_4_FBK,
      I2 => EXP5_EXP_PT_0_2_INV,
      I3 => EXP5_EXP_PT_0_3_INV,
      I4 => EXP5_EXP_PT_0_4_INV,
      I5 => EXP5_EXP_PT_0_5_INV,
      I6 => EXP5_EXP_PT_0_6_INV,
      I7 => EXP5_EXP_PT_0_7_INV,
      I8 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I9 => VCC,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP5_EXP_PT_0
    );
  EXP5_EXP_PT_1_639 : X_AND16 
    port map (
      I0 => EXP5_EXP_PT_1_0_INV,
      I1 => EXP5_EXP_PT_1_1_INV,
      I2 => EXP5_EXP_PT_1_2_INV,
      I3 => EXP5_EXP_PT_1_3_INV,
      I4 => EXP5_EXP_PT_1_4_INV,
      I5 => EXP5_EXP_PT_1_5_INV,
      I6 => EXP5_EXP_PT_1_6_INV,
      I7 => LIGHT_VALUE(5),
      I8 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I9 => VCC,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP5_EXP_PT_1
    );
  EXP5_EXP_PT_2_640 : X_AND16 
    port map (
      I0 => EXP5_EXP_PT_2_0_INV,
      I1 => EXP5_EXP_PT_2_1_INV,
      I2 => EXP5_EXP_PT_2_2_INV,
      I3 => EXP5_EXP_PT_2_3_INV,
      I4 => EXP5_EXP_PT_2_4_INV,
      I5 => EXP5_EXP_PT_2_5_INV,
      I6 => EXP5_EXP_PT_2_6_INV,
      I7 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      I8 => LIGHT_VALUE(0),
      I9 => VCC,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP5_EXP_PT_2
    );
  EXP5_EXP_PT_3_641 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => EXP5_EXP_PT_3_1_INV,
      I2 => FC1_CNT_3_FBK,
      I3 => FC1_CNT(1),
      I4 => FC1_CNT(2),
      I5 => FC1_CNT_4_FBK,
      I6 => FC1_CNT_5_FBK,
      I7 => FC1_CNT(0),
      I8 => EXP5_EXP_PT_3_8_INV,
      I9 => EXP5_EXP_PT_3_9_INV,
      I10 => VCC,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP5_EXP_PT_3
    );
  EXP5_EXP_PT_4_642 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      I1 => EXP5_EXP_PT_4_1_INV,
      I2 => FC1_CNT_3_FBK,
      I3 => FC1_CNT(1),
      I4 => FC1_CNT(2),
      I5 => FC1_CNT_4_FBK,
      I6 => FC1_CNT_5_FBK,
      I7 => FC1_CNT(0),
      I8 => EXP5_EXP_PT_4_8_INV,
      I9 => EXP5_EXP_PT_4_9_INV,
      I10 => EXP5_EXP_PT_4_10_INV,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => EXP5_EXP_PT_4
    );
  EXP5_EXP_643 : X_OR5 
    port map (
      I0 => EXP5_EXP_PT_0,
      I1 => EXP5_EXP_PT_1,
      I2 => EXP5_EXP_PT_2,
      I3 => EXP5_EXP_PT_3,
      I4 => EXP5_EXP_PT_4,
      O => EXP5_EXP
    );
  LIGHT_VALUE_0_Q_644 : X_BUF 
    port map (
      I => LIGHT_VALUE_0_Q,
      O => LIGHT_VALUE(0)
    );
  LIGHT_VALUE_0_R_OR_PRLD_645 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_0_RSTF,
      I1 => PRLD,
      O => LIGHT_VALUE_0_R_OR_PRLD
    );
  LIGHT_VALUE_0_REG : X_FF 
    port map (
      I => LIGHT_VALUE_0_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => LIGHT_VALUE_0_R_OR_PRLD,
      O => LIGHT_VALUE_0_Q
    );
  LIGHT_VALUE_0_RSTF_PT_0_646 : X_AND2 
    port map (
      I0 => LIGHT_VALUE_0_RSTF_PT_0_0_INV,
      I1 => LIGHT_VALUE_0_RSTF_PT_0_1_INV,
      O => LIGHT_VALUE_0_RSTF_PT_0
    );
  LIGHT_VALUE_0_RSTF_647 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_0_RSTF_PT_0,
      I1 => LIGHT_VALUE_0_RSTF_PT_0,
      O => LIGHT_VALUE_0_RSTF
    );
  LIGHT_VALUE_0_D1_648 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => LIGHT_VALUE_0_D1
    );
  LIGHT_VALUE_0_D2_PT_0_649 : X_AND2 
    port map (
      I0 => FC1_CNT_2_EXP,
      I1 => FC1_CNT_2_EXP,
      O => LIGHT_VALUE_0_D2_PT_0
    );
  LIGHT_VALUE_0_D2_PT_1_650 : X_AND2 
    port map (
      I0 => TD1_CNT_5_EXP,
      I1 => TD1_CNT_5_EXP,
      O => LIGHT_VALUE_0_D2_PT_1
    );
  LIGHT_VALUE_0_D2_PT_2_651 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => LIGHT_VALUE_0_D2_PT_2_1_INV,
      I2 => LIGHT_VALUE_0_D2_PT_2_2_INV,
      I3 => LIGHT_VALUE_0_D2_PT_2_3_INV,
      I4 => LIGHT_VALUE_0_D2_PT_2_4_INV,
      I5 => LIGHT_VALUE_0_D2_PT_2_5_INV,
      I6 => LIGHT_VALUE_0_D2_PT_2_6_INV,
      I7 => LIGHT_VALUE_0_D2_PT_2_7_INV,
      I8 => LIGHT_VALUE_0_D2_PT_2_8_INV,
      I9 => LIGHT_VALUE_0_D2_PT_2_9_INV,
      I10 => LIGHT_VALUE_1_FBK,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_0_D2_PT_2
    );
  LIGHT_VALUE_0_D2_PT_3_652 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => LIGHT_VALUE_0_D2_PT_3_1_INV,
      I2 => LIGHT_VALUE_0_D2_PT_3_2_INV,
      I3 => LIGHT_VALUE_0_D2_PT_3_3_INV,
      I4 => LIGHT_VALUE_0_D2_PT_3_4_INV,
      I5 => LIGHT_VALUE_0_D2_PT_3_5_INV,
      I6 => LIGHT_VALUE_0_D2_PT_3_6_INV,
      I7 => LIGHT_VALUE_0_D2_PT_3_7_INV,
      I8 => LIGHT_VALUE_0_D2_PT_3_8_INV,
      I9 => LIGHT_VALUE_0_D2_PT_3_9_INV,
      I10 => LIGHT_VALUE_2_FBK,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_0_D2_PT_3
    );
  LIGHT_VALUE_0_D2_PT_4_653 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => LIGHT_VALUE_0_D2_PT_4_1_INV,
      I2 => LIGHT_VALUE_0_D2_PT_4_2_INV,
      I3 => LIGHT_VALUE_0_D2_PT_4_3_INV,
      I4 => LIGHT_VALUE_0_D2_PT_4_4_INV,
      I5 => LIGHT_VALUE_0_D2_PT_4_5_INV,
      I6 => LIGHT_VALUE_0_D2_PT_4_6_INV,
      I7 => LIGHT_VALUE_0_D2_PT_4_7_INV,
      I8 => LIGHT_VALUE_0_D2_PT_4_8_INV,
      I9 => LIGHT_VALUE_0_D2_PT_4_9_INV,
      I10 => LIGHT_VALUE_3_FBK,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_0_D2_PT_4
    );
  LIGHT_VALUE_0_D2_PT_5_654 : X_AND16 
    port map (
      I0 => LIGHT_VALUE_0_D2_PT_5_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I2 => LIGHT_VALUE_0_D2_PT_5_2_INV,
      I3 => FC1_CNT_1_FBK,
      I4 => FC1_CNT_2_FBK,
      I5 => FC1_CNT_0_FBK,
      I6 => FC1_CNT(3),
      I7 => FC1_CNT(4),
      I8 => FC1_CNT(5),
      I9 => FC1_CNT(6),
      I10 => FC1_CNT(7),
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_0_D2_PT_5
    );
  LIGHT_VALUE_0_D2_655 : X_OR6 
    port map (
      I0 => LIGHT_VALUE_0_D2_PT_0,
      I1 => LIGHT_VALUE_0_D2_PT_1,
      I2 => LIGHT_VALUE_0_D2_PT_2,
      I3 => LIGHT_VALUE_0_D2_PT_3,
      I4 => LIGHT_VALUE_0_D2_PT_4,
      I5 => LIGHT_VALUE_0_D2_PT_5,
      O => LIGHT_VALUE_0_D2
    );
  LIGHT_VALUE_0_D_656 : X_XOR2 
    port map (
      I0 => LIGHT_VALUE_0_D_TFF,
      I1 => LIGHT_VALUE_0_Q,
      O => LIGHT_VALUE_0_D
    );
  LIGHT_VALUE_0_XOR : X_XOR2 
    port map (
      I0 => LIGHT_VALUE_0_D1,
      I1 => LIGHT_VALUE_0_D2,
      O => LIGHT_VALUE_0_D_TFF
    );
  LIGHT_VALUE_0_FBK_657 : X_BUF 
    port map (
      I => LIGHT_VALUE_0_Q,
      O => LIGHT_VALUE_0_FBK
    );
  TD1_CNT_5_Q_658 : X_BUF 
    port map (
      I => TD1_CNT_5_Q,
      O => TD1_CNT_5_Q_0
    );
  TD1_CNT_5_REG : X_FF 
    port map (
      I => TD1_CNT_5_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => TD1_CNT_5_SETF,
      RST => PRLD,
      O => TD1_CNT_5_Q
    );
  TD1_CNT_5_SETF_PT_0_659 : X_AND2 
    port map (
      I0 => TD1_CNT_5_SETF_PT_0_0_INV,
      I1 => TD1_CNT_5_SETF_PT_0_1_INV,
      O => TD1_CNT_5_SETF_PT_0
    );
  TD1_CNT_5_SETF_660 : X_OR2 
    port map (
      I0 => TD1_CNT_5_SETF_PT_0,
      I1 => TD1_CNT_5_SETF_PT_0,
      O => TD1_CNT_5_SETF
    );
  TD1_CNT_5_D1_661 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => TD1_CNT_5_D1
    );
  TD1_CNT_5_D2_PT_0_662 : X_AND5 
    port map (
      I0 => TD1_CNT_5_D2_PT_0_0_INV,
      I1 => TD1_CNT_5_D2_PT_0_1_INV,
      I2 => TD1_CNT_5_D2_PT_0_2_INV,
      I3 => TD1_CNT_5_D2_PT_0_3_INV,
      I4 => TD1_CNT_5_D2_PT_0_4_INV,
      O => TD1_CNT_5_D2_PT_0
    );
  TD1_CNT_5_D2_663 : X_OR2 
    port map (
      I0 => TD1_CNT_5_D2_PT_0,
      I1 => TD1_CNT_5_D2_PT_0,
      O => TD1_CNT_5_D2
    );
  TD1_CNT_5_D_664 : X_XOR2 
    port map (
      I0 => TD1_CNT_5_D_TFF,
      I1 => TD1_CNT_5_Q,
      O => TD1_CNT_5_D
    );
  TD1_CNT_5_XOR : X_XOR2 
    port map (
      I0 => TD1_CNT_5_D1,
      I1 => TD1_CNT_5_D2,
      O => TD1_CNT_5_D_TFF
    );
  TD1_CNT_5_EXP_PT_0_665 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => TD1_CNT_5_EXP_PT_0_1_INV,
      I2 => LIGHT_VALUE_5_FBK,
      I3 => TD1_CNT_5_EXP_PT_0_3_INV,
      I4 => TD1_CNT_5_EXP_PT_0_4_INV,
      I5 => TD1_CNT_5_EXP_PT_0_5_INV,
      I6 => TD1_CNT_5_EXP_PT_0_6_INV,
      I7 => TD1_CNT_5_EXP_PT_0_7_INV,
      I8 => TD1_CNT_5_EXP_PT_0_8_INV,
      I9 => TD1_CNT_5_EXP_PT_0_9_INV,
      I10 => TD1_CNT_5_EXP_PT_0_10_INV,
      I11 => VCC,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => TD1_CNT_5_EXP_PT_0
    );
  TD1_CNT_5_EXP_PT_1_666 : X_AND16 
    port map (
      I0 => TD1_CNT_5_EXP_PT_1_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I2 => FC1_CNT_1_FBK,
      I3 => FC1_CNT_2_FBK,
      I4 => FC1_CNT_0_FBK,
      I5 => FC1_CNT(3),
      I6 => FC1_CNT(4),
      I7 => FC1_CNT(5),
      I8 => FC1_CNT(6),
      I9 => FC1_CNT(7),
      I10 => TD1_CNT_5_EXP_PT_1_10_INV,
      I11 => TD1_CNT_5_EXP_PT_1_11_INV,
      I12 => VCC,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => TD1_CNT_5_EXP_PT_1
    );
  TD1_CNT_5_EXP_PT_2_667 : X_AND16 
    port map (
      I0 => TD1_CNT_5_EXP_PT_2_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I2 => FC1_CNT_1_FBK,
      I3 => FC1_CNT_2_FBK,
      I4 => FC1_CNT_0_FBK,
      I5 => FC1_CNT(3),
      I6 => FC1_CNT(4),
      I7 => FC1_CNT(5),
      I8 => FC1_CNT(6),
      I9 => FC1_CNT(7),
      I10 => TD1_CNT_5_EXP_PT_2_10_INV,
      I11 => TD1_CNT_5_EXP_PT_2_11_INV,
      I12 => TD1_CNT_5_EXP_PT_2_12_INV,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => TD1_CNT_5_EXP_PT_2
    );
  TD1_CNT_5_EXP_668 : X_OR3 
    port map (
      I0 => TD1_CNT_5_EXP_PT_0,
      I1 => TD1_CNT_5_EXP_PT_1,
      I2 => TD1_CNT_5_EXP_PT_2,
      O => TD1_CNT_5_EXP
    );
  TD1_CNT_1_Q_669 : X_BUF 
    port map (
      I => TD1_CNT_1_Q,
      O => TD1_CNT_1_Q_3
    );
  TD1_CNT_1_REG : X_FF 
    port map (
      I => TD1_CNT_1_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => TD1_CNT_1_SETF,
      RST => PRLD,
      O => TD1_CNT_1_Q
    );
  TD1_CNT_1_SETF_PT_0_670 : X_AND2 
    port map (
      I0 => TD1_CNT_1_SETF_PT_0_0_INV,
      I1 => TD1_CNT_1_SETF_PT_0_1_INV,
      O => TD1_CNT_1_SETF_PT_0
    );
  TD1_CNT_1_SETF_671 : X_OR2 
    port map (
      I0 => TD1_CNT_1_SETF_PT_0,
      I1 => TD1_CNT_1_SETF_PT_0,
      O => TD1_CNT_1_SETF
    );
  TD1_CNT_1_D1_672 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => TD1_CNT_1_D1
    );
  TD1_CNT_1_D2_PT_0_673 : X_AND2 
    port map (
      I0 => TD1_CNT_0_Q_2,
      I1 => TD1_CNT_0_Q_2,
      O => TD1_CNT_1_D2_PT_0
    );
  TD1_CNT_1_D2_674 : X_OR2 
    port map (
      I0 => TD1_CNT_1_D2_PT_0,
      I1 => TD1_CNT_1_D2_PT_0,
      O => TD1_CNT_1_D2
    );
  TD1_CNT_1_D_675 : X_XOR2 
    port map (
      I0 => TD1_CNT_1_D_TFF,
      I1 => TD1_CNT_1_Q,
      O => TD1_CNT_1_D
    );
  TD1_CNT_1_XOR : X_XOR2 
    port map (
      I0 => TD1_CNT_1_XOR_0_INV,
      I1 => TD1_CNT_1_D2,
      O => TD1_CNT_1_D_TFF
    );
  TD1_CNT_2_FBK_676 : X_BUF 
    port map (
      I => TD1_CNT_2_Q,
      O => TD1_CNT_2_FBK
    );
  TD1_CNT_2_R_OR_PRLD_677 : X_OR2 
    port map (
      I0 => TD1_CNT_2_RSTF,
      I1 => PRLD,
      O => TD1_CNT_2_R_OR_PRLD
    );
  TD1_CNT_2_REG : X_FF 
    port map (
      I => TD1_CNT_2_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => TD1_CNT_2_R_OR_PRLD,
      O => TD1_CNT_2_Q
    );
  TD1_CNT_2_RSTF_PT_0_678 : X_AND2 
    port map (
      I0 => TD1_CNT_2_RSTF_PT_0_0_INV,
      I1 => TD1_CNT_2_RSTF_PT_0_1_INV,
      O => TD1_CNT_2_RSTF_PT_0
    );
  TD1_CNT_2_RSTF_679 : X_OR2 
    port map (
      I0 => TD1_CNT_2_RSTF_PT_0,
      I1 => TD1_CNT_2_RSTF_PT_0,
      O => TD1_CNT_2_RSTF
    );
  TD1_CNT_2_D1_680 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => TD1_CNT_2_D1
    );
  TD1_CNT_2_D2_PT_0_681 : X_AND2 
    port map (
      I0 => TD1_CNT_2_D2_PT_0_0_INV,
      I1 => TD1_CNT_2_D2_PT_0_1_INV,
      O => TD1_CNT_2_D2_PT_0
    );
  TD1_CNT_2_D2_682 : X_OR2 
    port map (
      I0 => TD1_CNT_2_D2_PT_0,
      I1 => TD1_CNT_2_D2_PT_0,
      O => TD1_CNT_2_D2
    );
  TD1_CNT_2_D_683 : X_XOR2 
    port map (
      I0 => TD1_CNT_2_D_TFF,
      I1 => TD1_CNT_2_Q,
      O => TD1_CNT_2_D
    );
  TD1_CNT_2_XOR : X_XOR2 
    port map (
      I0 => TD1_CNT_2_D1,
      I1 => TD1_CNT_2_D2,
      O => TD1_CNT_2_D_TFF
    );
  TD1_CNT_3_EXP_PT_0_684 : X_AND5 
    port map (
      I0 => TD1_CNT_3_EXP_PT_0_0_INV,
      I1 => TD1_CNT_3_EXP_PT_0_1_INV,
      I2 => TD1_CNT_3_EXP_PT_0_2_INV,
      I3 => TD1_CNT_3_EXP_PT_0_3_INV,
      I4 => TD1_CNT_0_FBK,
      O => TD1_CNT_3_EXP_PT_0
    );
  TD1_CNT_3_EXP_PT_1_685 : X_AND5 
    port map (
      I0 => TD1_CNT_3_EXP_PT_1_0_INV,
      I1 => TD1_CNT_3_EXP_PT_1_1_INV,
      I2 => TD1_CNT_3_EXP_PT_1_2_INV,
      I3 => TD1_CNT_0_FBK,
      I4 => TD1_CNT_1_Q_3,
      O => TD1_CNT_3_EXP_PT_1
    );
  TD1_CNT_3_EXP_686 : X_OR2 
    port map (
      I0 => TD1_CNT_3_EXP_PT_0,
      I1 => TD1_CNT_3_EXP_PT_1,
      O => TD1_CNT_3_EXP
    );
  TD1_CNT_3_FBK_687 : X_BUF 
    port map (
      I => TD1_CNT_3_Q,
      O => TD1_CNT_3_FBK
    );
  TD1_CNT_3_REG : X_FF 
    port map (
      I => TD1_CNT_3_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => TD1_CNT_3_SETF,
      RST => PRLD,
      O => TD1_CNT_3_Q
    );
  TD1_CNT_3_SETF_PT_0_688 : X_AND2 
    port map (
      I0 => TD1_CNT_3_SETF_PT_0_0_INV,
      I1 => TD1_CNT_3_SETF_PT_0_1_INV,
      O => TD1_CNT_3_SETF_PT_0
    );
  TD1_CNT_3_SETF_689 : X_OR2 
    port map (
      I0 => TD1_CNT_3_SETF_PT_0,
      I1 => TD1_CNT_3_SETF_PT_0,
      O => TD1_CNT_3_SETF
    );
  TD1_CNT_3_D1_690 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => TD1_CNT_3_D1
    );
  TD1_CNT_3_D2_PT_0_691 : X_AND3 
    port map (
      I0 => TD1_CNT_3_D2_PT_0_0_INV,
      I1 => TD1_CNT_3_D2_PT_0_1_INV,
      I2 => TD1_CNT_3_D2_PT_0_2_INV,
      O => TD1_CNT_3_D2_PT_0
    );
  TD1_CNT_3_D2_692 : X_OR2 
    port map (
      I0 => TD1_CNT_3_D2_PT_0,
      I1 => TD1_CNT_3_D2_PT_0,
      O => TD1_CNT_3_D2
    );
  TD1_CNT_3_D_693 : X_XOR2 
    port map (
      I0 => TD1_CNT_3_D_TFF,
      I1 => TD1_CNT_3_Q,
      O => TD1_CNT_3_D
    );
  TD1_CNT_3_XOR : X_XOR2 
    port map (
      I0 => TD1_CNT_3_D1,
      I1 => TD1_CNT_3_D2,
      O => TD1_CNT_3_D_TFF
    );
  LIGHT_VALUE_2_Q_694 : X_BUF 
    port map (
      I => LIGHT_VALUE_2_Q,
      O => LIGHT_VALUE(2)
    );
  LIGHT_VALUE_2_R_OR_PRLD_695 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_2_RSTF,
      I1 => PRLD,
      O => LIGHT_VALUE_2_R_OR_PRLD
    );
  LIGHT_VALUE_2_REG : X_FF 
    port map (
      I => LIGHT_VALUE_2_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => LIGHT_VALUE_2_R_OR_PRLD,
      O => LIGHT_VALUE_2_Q
    );
  LIGHT_VALUE_2_RSTF_PT_0_696 : X_AND2 
    port map (
      I0 => LIGHT_VALUE_2_RSTF_PT_0_0_INV,
      I1 => LIGHT_VALUE_2_RSTF_PT_0_1_INV,
      O => LIGHT_VALUE_2_RSTF_PT_0
    );
  LIGHT_VALUE_2_RSTF_697 : X_OR2 
    port map (
      I0 => LIGHT_VALUE_2_RSTF_PT_0,
      I1 => LIGHT_VALUE_2_RSTF_PT_0,
      O => LIGHT_VALUE_2_RSTF
    );
  LIGHT_VALUE_2_D1_698 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => LIGHT_VALUE_2_D1
    );
  LIGHT_VALUE_2_D2_PT_0_699 : X_AND2 
    port map (
      I0 => LIGHT_VALUE_3_EXP,
      I1 => LIGHT_VALUE_3_EXP,
      O => LIGHT_VALUE_2_D2_PT_0
    );
  LIGHT_VALUE_2_D2_PT_1_700 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => LIGHT_VALUE_2_D2_PT_1_1_INV,
      I2 => LIGHT_VALUE_2_D2_PT_1_2_INV,
      I3 => LIGHT_VALUE_2_D2_PT_1_3_INV,
      I4 => LIGHT_VALUE_2_D2_PT_1_4_INV,
      I5 => LIGHT_VALUE_2_D2_PT_1_5_INV,
      I6 => LIGHT_VALUE_2_D2_PT_1_6_INV,
      I7 => LIGHT_VALUE_2_D2_PT_1_7_INV,
      I8 => LIGHT_VALUE_2_D2_PT_1_8_INV,
      I9 => LIGHT_VALUE_2_D2_PT_1_9_INV,
      I10 => LIGHT_VALUE_2_D2_PT_1_10_INV,
      I11 => LIGHT_VALUE_2_FBK,
      I12 => LIGHT_VALUE_2_D2_PT_1_12_INV,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_2_D2_PT_1
    );
  LIGHT_VALUE_2_D2_PT_2_701 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => LIGHT_VALUE_2_D2_PT_2_1_INV,
      I2 => LIGHT_VALUE_2_D2_PT_2_2_INV,
      I3 => LIGHT_VALUE_2_D2_PT_2_3_INV,
      I4 => LIGHT_VALUE_2_D2_PT_2_4_INV,
      I5 => LIGHT_VALUE_2_D2_PT_2_5_INV,
      I6 => LIGHT_VALUE_2_D2_PT_2_6_INV,
      I7 => LIGHT_VALUE_2_D2_PT_2_7_INV,
      I8 => LIGHT_VALUE_2_D2_PT_2_8_INV,
      I9 => LIGHT_VALUE_2_D2_PT_2_9_INV,
      I10 => LIGHT_VALUE_2_D2_PT_2_10_INV,
      I11 => LIGHT_VALUE_2_D2_PT_2_11_INV,
      I12 => LIGHT_VALUE_3_FBK,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_2_D2_PT_2
    );
  LIGHT_VALUE_2_D2_PT_3_702 : X_AND16 
    port map (
      I0 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      I1 => LIGHT_VALUE_2_D2_PT_3_1_INV,
      I2 => LIGHT_VALUE_2_D2_PT_3_2_INV,
      I3 => LIGHT_VALUE_2_D2_PT_3_3_INV,
      I4 => LIGHT_VALUE_2_D2_PT_3_4_INV,
      I5 => LIGHT_VALUE_2_D2_PT_3_5_INV,
      I6 => LIGHT_VALUE_2_D2_PT_3_6_INV,
      I7 => LIGHT_VALUE_2_D2_PT_3_7_INV,
      I8 => LIGHT_VALUE_2_D2_PT_3_8_INV,
      I9 => LIGHT_VALUE_2_D2_PT_3_9_INV,
      I10 => LIGHT_VALUE_2_D2_PT_3_10_INV,
      I11 => LIGHT_VALUE_2_D2_PT_3_11_INV,
      I12 => LIGHT_VALUE(4),
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_2_D2_PT_3
    );
  LIGHT_VALUE_2_D2_PT_4_703 : X_AND16 
    port map (
      I0 => LIGHT_VALUE_2_D2_PT_4_0_INV,
      I1 => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      I2 => LIGHT_VALUE_2_D2_PT_4_2_INV,
      I3 => FC1_CNT_1_FBK,
      I4 => FC1_CNT_2_FBK,
      I5 => FC1_CNT_0_FBK,
      I6 => FC1_CNT(3),
      I7 => FC1_CNT(4),
      I8 => FC1_CNT(5),
      I9 => FC1_CNT(6),
      I10 => FC1_CNT(7),
      I11 => LIGHT_VALUE_1_FBK,
      I12 => LIGHT_VALUE_0_FBK,
      I13 => VCC,
      I14 => VCC,
      I15 => VCC,
      O => LIGHT_VALUE_2_D2_PT_4
    );
  LIGHT_VALUE_2_D2_704 : X_OR5 
    port map (
      I0 => LIGHT_VALUE_2_D2_PT_0,
      I1 => LIGHT_VALUE_2_D2_PT_1,
      I2 => LIGHT_VALUE_2_D2_PT_2,
      I3 => LIGHT_VALUE_2_D2_PT_3,
      I4 => LIGHT_VALUE_2_D2_PT_4,
      O => LIGHT_VALUE_2_D2
    );
  LIGHT_VALUE_2_D_705 : X_XOR2 
    port map (
      I0 => LIGHT_VALUE_2_D_TFF,
      I1 => LIGHT_VALUE_2_Q,
      O => LIGHT_VALUE_2_D
    );
  LIGHT_VALUE_2_XOR : X_XOR2 
    port map (
      I0 => LIGHT_VALUE_2_D1,
      I1 => LIGHT_VALUE_2_D2,
      O => LIGHT_VALUE_2_D_TFF
    );
  LIGHT_VALUE_2_FBK_706 : X_BUF 
    port map (
      I => LIGHT_VALUE_2_Q,
      O => LIGHT_VALUE_2_FBK
    );
  TD1_CNT_4_Q_707 : X_BUF 
    port map (
      I => TD1_CNT_4_Q,
      O => TD1_CNT_4_Q_1
    );
  TD1_CNT_4_R_OR_PRLD_708 : X_OR2 
    port map (
      I0 => TD1_CNT_4_RSTF,
      I1 => PRLD,
      O => TD1_CNT_4_R_OR_PRLD
    );
  TD1_CNT_4_REG : X_FF 
    port map (
      I => TD1_CNT_4_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => TD1_CNT_4_R_OR_PRLD,
      O => TD1_CNT_4_Q
    );
  TD1_CNT_4_RSTF_PT_0_709 : X_AND2 
    port map (
      I0 => TD1_CNT_4_RSTF_PT_0_0_INV,
      I1 => TD1_CNT_4_RSTF_PT_0_1_INV,
      O => TD1_CNT_4_RSTF_PT_0
    );
  TD1_CNT_4_RSTF_710 : X_OR2 
    port map (
      I0 => TD1_CNT_4_RSTF_PT_0,
      I1 => TD1_CNT_4_RSTF_PT_0,
      O => TD1_CNT_4_RSTF
    );
  TD1_CNT_4_D1_711 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => TD1_CNT_4_D1
    );
  TD1_CNT_4_D2_PT_0_712 : X_AND4 
    port map (
      I0 => TD1_CNT_4_D2_PT_0_0_INV,
      I1 => TD1_CNT_4_D2_PT_0_1_INV,
      I2 => TD1_CNT_4_D2_PT_0_2_INV,
      I3 => TD1_CNT_4_D2_PT_0_3_INV,
      O => TD1_CNT_4_D2_PT_0
    );
  TD1_CNT_4_D2_713 : X_OR2 
    port map (
      I0 => TD1_CNT_4_D2_PT_0,
      I1 => TD1_CNT_4_D2_PT_0,
      O => TD1_CNT_4_D2
    );
  TD1_CNT_4_D_714 : X_XOR2 
    port map (
      I0 => TD1_CNT_4_D_TFF,
      I1 => TD1_CNT_4_Q,
      O => TD1_CNT_4_D
    );
  TD1_CNT_4_XOR : X_XOR2 
    port map (
      I0 => TD1_CNT_4_D1,
      I1 => TD1_CNT_4_D2,
      O => TD1_CNT_4_D_TFF
    );
  TD1_CNT_4_EXP_PT_0_715 : X_AND4 
    port map (
      I0 => TD1_CNT_4_EXP_PT_0_0_INV,
      I1 => TD1_CNT_4_EXP_PT_0_1_INV,
      I2 => TD1_CNT_4_EXP_PT_0_2_INV,
      I3 => TD1_CNT_1_Q_3,
      O => TD1_CNT_4_EXP_PT_0
    );
  TD1_CNT_4_EXP_PT_1_716 : X_AND4 
    port map (
      I0 => TD1_CNT_4_EXP_PT_1_0_INV,
      I1 => TD1_CNT_4_EXP_PT_1_1_INV,
      I2 => TD1_CNT_1_Q_3,
      I3 => TD1_CNT_2_FBK,
      O => TD1_CNT_4_EXP_PT_1
    );
  TD1_CNT_4_EXP_PT_2_717 : X_AND5 
    port map (
      I0 => TD1_CNT_4_EXP_PT_2_0_INV,
      I1 => TD1_CNT_0_FBK,
      I2 => TD1_CNT_1_Q_3,
      I3 => TD1_CNT_2_FBK,
      I4 => TD1_CNT_3_FBK,
      O => TD1_CNT_4_EXP_PT_2
    );
  TD1_CNT_4_EXP_718 : X_OR3 
    port map (
      I0 => TD1_CNT_4_EXP_PT_0,
      I1 => TD1_CNT_4_EXP_PT_1,
      I2 => TD1_CNT_4_EXP_PT_2,
      O => TD1_CNT_4_EXP
    );
  TD1_CNT_4_FBK_719 : X_BUF 
    port map (
      I => TD1_CNT_4_Q,
      O => TD1_CNT_4_FBK
    );
  CM_FADE_UP_720 : X_BUF 
    port map (
      I => CM_FADE_UP_Q,
      O => CM_FADE_UP
    );
  CM_FADE_UP_R_OR_PRLD_721 : X_OR2 
    port map (
      I0 => FSRIO_0,
      I1 => PRLD,
      O => CM_FADE_UP_R_OR_PRLD
    );
  CM_FADE_UP_REG : X_FF 
    port map (
      I => CM_FADE_UP_D,
      CLK => CLK_C_FCLK,
      CE => VCC,
      SET => GND,
      RST => CM_FADE_UP_R_OR_PRLD,
      O => CM_FADE_UP_Q
    );
  CM_FADE_UP_D1_722 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => CM_FADE_UP_D1
    );
  CM_FADE_UP_D2_PT_0_723 : X_AND2 
    port map (
      I0 => RXD_ACK,
      I1 => RXD_ACK,
      O => CM_FADE_UP_D2_PT_0
    );
  CM_FADE_UP_D2_PT_1_724 : X_AND2 
    port map (
      I0 => RXD_2_FBK,
      I1 => RXD_2_FBK,
      O => CM_FADE_UP_D2_PT_1
    );
  CM_FADE_UP_D2_PT_2_725 : X_AND2 
    port map (
      I0 => CM_FADE_UP_D2_PT_2_0_INV,
      I1 => CM_FADE_UP_D2_PT_2_1_INV,
      O => CM_FADE_UP_D2_PT_2
    );
  CM_FADE_UP_D2_PT_3_726 : X_AND2 
    port map (
      I0 => EXP15_EXP,
      I1 => EXP15_EXP,
      O => CM_FADE_UP_D2_PT_3
    );
  CM_FADE_UP_D2_PT_4_727 : X_AND2 
    port map (
      I0 => RXD_READY_EXP,
      I1 => RXD_READY_EXP,
      O => CM_FADE_UP_D2_PT_4
    );
  CM_FADE_UP_D2_PT_5_728 : X_AND2 
    port map (
      I0 => RC_ADDRESS_C(0),
      I1 => CM_FADE_UP_D2_PT_5_1_INV,
      O => CM_FADE_UP_D2_PT_5
    );
  CM_FADE_UP_D2_PT_6_729 : X_AND2 
    port map (
      I0 => CM_FADE_UP_D2_PT_6_0_INV,
      I1 => RXD_4_FBK,
      O => CM_FADE_UP_D2_PT_6
    );
  CM_FADE_UP_D2_730 : X_OR7 
    port map (
      I0 => CM_FADE_UP_D2_PT_0,
      I1 => CM_FADE_UP_D2_PT_1,
      I2 => CM_FADE_UP_D2_PT_2,
      I3 => CM_FADE_UP_D2_PT_3,
      I4 => CM_FADE_UP_D2_PT_4,
      I5 => CM_FADE_UP_D2_PT_5,
      I6 => CM_FADE_UP_D2_PT_6,
      O => CM_FADE_UP_D2
    );
  CM_FADE_UP_D_731 : X_XOR2 
    port map (
      I0 => CM_FADE_UP_D_TFF,
      I1 => CM_FADE_UP_Q,
      O => CM_FADE_UP_D
    );
  CM_FADE_UP_XOR : X_XOR2 
    port map (
      I0 => CM_FADE_UP_XOR_0_INV,
      I1 => CM_FADE_UP_D2,
      O => CM_FADE_UP_D_TFF
    );
  CM_FADE_UP_FBK_732 : X_BUF 
    port map (
      I => CM_FADE_UP_Q,
      O => CM_FADE_UP_FBK
    );
  EXP15_EXP_PT_0_733 : X_AND2 
    port map (
      I0 => EXP16_EXP,
      I1 => EXP16_EXP,
      O => EXP15_EXP_PT_0
    );
  EXP15_EXP_PT_1_734 : X_AND2 
    port map (
      I0 => RXD_3_FBK,
      I1 => EXP15_EXP_PT_1_1_INV,
      O => EXP15_EXP_PT_1
    );
  EXP15_EXP_PT_2_735 : X_AND2 
    port map (
      I0 => RXD_1_FBK,
      I1 => CM_FADE_UP_FBK,
      O => EXP15_EXP_PT_2
    );
  EXP15_EXP_PT_3_736 : X_AND2 
    port map (
      I0 => EXP15_EXP_PT_3_0_INV,
      I1 => EXP15_EXP_PT_3_1_INV,
      O => EXP15_EXP_PT_3
    );
  EXP15_EXP_PT_4_737 : X_AND2 
    port map (
      I0 => RXD_0_FBK,
      I1 => EXP15_EXP_PT_4_1_INV,
      O => EXP15_EXP_PT_4
    );
  EXP15_EXP_PT_5_738 : X_AND2 
    port map (
      I0 => EXP15_EXP_PT_5_0_INV,
      I1 => RXD_7_FBK,
      O => EXP15_EXP_PT_5
    );
  EXP15_EXP_739 : X_OR6 
    port map (
      I0 => EXP15_EXP_PT_0,
      I1 => EXP15_EXP_PT_1,
      I2 => EXP15_EXP_PT_2,
      I3 => EXP15_EXP_PT_3,
      I4 => EXP15_EXP_PT_4,
      I5 => EXP15_EXP_PT_5,
      O => EXP15_EXP
    );
  EXP16_EXP_PT_0_740 : X_AND2 
    port map (
      I0 => RXD_3_FBK,
      I1 => RXD_0_FBK,
      O => EXP16_EXP_PT_0
    );
  EXP16_EXP_PT_1_741 : X_AND3 
    port map (
      I0 => EXP16_EXP_PT_1_0_INV,
      I1 => EXP16_EXP_PT_1_1_INV,
      I2 => CM_FADE_UP_FBK,
      O => EXP16_EXP_PT_1
    );
  EXP16_EXP_742 : X_OR2 
    port map (
      I0 => EXP16_EXP_PT_0,
      I1 => EXP16_EXP_PT_1,
      O => EXP16_EXP
    );
  Q_OPTX_FX_DC_68_UIM_743 : X_BUF 
    port map (
      I => Q_OPTX_FX_DC_68_Q,
      O => Q_OPTX_FX_DC_68_UIM
    );
  Q_OPTX_FX_DC_68_REG : X_BUF 
    port map (
      I => Q_OPTX_FX_DC_68_D,
      O => Q_OPTX_FX_DC_68_Q
    );
  Q_OPTX_FX_DC_68_D1_744 : X_OR2 
    port map (
      I0 => GND,
      I1 => GND,
      O => Q_OPTX_FX_DC_68_D1
    );
  Q_OPTX_FX_DC_68_D2_PT_0_745 : X_AND2 
    port map (
      I0 => TD1_CNT_4_EXP,
      I1 => TD1_CNT_4_EXP,
      O => Q_OPTX_FX_DC_68_D2_PT_0
    );
  Q_OPTX_FX_DC_68_D2_PT_1_746 : X_AND2 
    port map (
      I0 => EXP11_EXP,
      I1 => EXP11_EXP,
      O => Q_OPTX_FX_DC_68_D2_PT_1
    );
  Q_OPTX_FX_DC_68_D2_PT_2_747 : X_AND2 
    port map (
      I0 => Q_OPTX_FX_DC_68_D2_PT_2_0_INV,
      I1 => TD1_CNT_3_FBK,
      O => Q_OPTX_FX_DC_68_D2_PT_2
    );
  Q_OPTX_FX_DC_68_D2_PT_3_748 : X_AND3 
    port map (
      I0 => Q_OPTX_FX_DC_68_D2_PT_3_0_INV,
      I1 => Q_OPTX_FX_DC_68_D2_PT_3_1_INV,
      I2 => TD1_CNT_2_FBK,
      O => Q_OPTX_FX_DC_68_D2_PT_3
    );
  Q_OPTX_FX_DC_68_D2_PT_4_749 : X_AND3 
    port map (
      I0 => Q_OPTX_FX_DC_68_D2_PT_4_0_INV,
      I1 => TD1_CNT_2_FBK,
      I2 => TD1_CNT_3_FBK,
      O => Q_OPTX_FX_DC_68_D2_PT_4
    );
  Q_OPTX_FX_DC_68_D2_PT_5_750 : X_AND4 
    port map (
      I0 => Q_OPTX_FX_DC_68_D2_PT_5_0_INV,
      I1 => Q_OPTX_FX_DC_68_D2_PT_5_1_INV,
      I2 => TD1_CNT_1_Q_3,
      I3 => TD1_CNT_3_FBK,
      O => Q_OPTX_FX_DC_68_D2_PT_5
    );
  Q_OPTX_FX_DC_68_D2_PT_6_751 : X_AND4 
    port map (
      I0 => Q_OPTX_FX_DC_68_D2_PT_6_0_INV,
      I1 => TD1_CNT_1_Q_3,
      I2 => TD1_CNT_2_FBK,
      I3 => TD1_CNT_3_FBK,
      O => Q_OPTX_FX_DC_68_D2_PT_6
    );
  Q_OPTX_FX_DC_68_D2_752 : X_OR7 
    port map (
      I0 => Q_OPTX_FX_DC_68_D2_PT_0,
      I1 => Q_OPTX_FX_DC_68_D2_PT_1,
      I2 => Q_OPTX_FX_DC_68_D2_PT_2,
      I3 => Q_OPTX_FX_DC_68_D2_PT_3,
      I4 => Q_OPTX_FX_DC_68_D2_PT_4,
      I5 => Q_OPTX_FX_DC_68_D2_PT_5,
      I6 => Q_OPTX_FX_DC_68_D2_PT_6,
      O => Q_OPTX_FX_DC_68_D2
    );
  Q_OPTX_FX_DC_68_XOR : X_XOR2 
    port map (
      I0 => Q_OPTX_FX_DC_68_D1,
      I1 => Q_OPTX_FX_DC_68_D2,
      O => Q_OPTX_FX_DC_68_D
    );
  EXP11_EXP_PT_0_753 : X_AND2 
    port map (
      I0 => TD1_CNT_3_EXP,
      I1 => TD1_CNT_3_EXP,
      O => EXP11_EXP_PT_0
    );
  EXP11_EXP_PT_1_754 : X_AND5 
    port map (
      I0 => EXP11_EXP_PT_1_0_INV,
      I1 => EXP11_EXP_PT_1_1_INV,
      I2 => EXP11_EXP_PT_1_2_INV,
      I3 => TD1_CNT_0_FBK,
      I4 => TD1_CNT_3_FBK,
      O => EXP11_EXP_PT_1
    );
  EXP11_EXP_PT_2_755 : X_AND5 
    port map (
      I0 => EXP11_EXP_PT_2_0_INV,
      I1 => EXP11_EXP_PT_2_1_INV,
      I2 => EXP11_EXP_PT_2_2_INV,
      I3 => TD1_CNT_0_FBK,
      I4 => TD1_CNT_2_FBK,
      O => EXP11_EXP_PT_2
    );
  EXP11_EXP_PT_3_756 : X_AND5 
    port map (
      I0 => EXP11_EXP_PT_3_0_INV,
      I1 => EXP11_EXP_PT_3_1_INV,
      I2 => TD1_CNT_0_FBK,
      I3 => TD1_CNT_2_FBK,
      I4 => TD1_CNT_3_FBK,
      O => EXP11_EXP_PT_3
    );
  EXP11_EXP_PT_4_757 : X_AND5 
    port map (
      I0 => EXP11_EXP_PT_4_0_INV,
      I1 => EXP11_EXP_PT_4_1_INV,
      I2 => TD1_CNT_0_FBK,
      I3 => TD1_CNT_1_Q_3,
      I4 => TD1_CNT_3_FBK,
      O => EXP11_EXP_PT_4
    );
  EXP11_EXP_PT_5_758 : X_AND5 
    port map (
      I0 => EXP11_EXP_PT_5_0_INV,
      I1 => EXP11_EXP_PT_5_1_INV,
      I2 => TD1_CNT_0_FBK,
      I3 => TD1_CNT_1_Q_3,
      I4 => TD1_CNT_2_FBK,
      O => EXP11_EXP_PT_5
    );
  EXP11_EXP_759 : X_OR6 
    port map (
      I0 => EXP11_EXP_PT_0,
      I1 => EXP11_EXP_PT_1,
      I2 => EXP11_EXP_PT_2,
      I3 => EXP11_EXP_PT_3,
      I4 => EXP11_EXP_PT_4,
      I5 => EXP11_EXP_PT_5,
      O => EXP11_EXP
    );
  TD1_TRIAC_TRIG_I_D2_PT_1_0_INV_760 : X_INV 
    port map (
      I => LIGHT_VALUE(5),
      O => TD1_TRIAC_TRIG_I_D2_PT_1_0_INV
    );
  TD1_TRIAC_TRIG_I_D2_PT_2_0_INV_761 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => TD1_TRIAC_TRIG_I_D2_PT_2_0_INV
    );
  TD1_TRIAC_TRIG_I_D2_PT_2_1_INV_762 : X_INV 
    port map (
      I => LIGHT_VALUE(5),
      O => TD1_TRIAC_TRIG_I_D2_PT_2_1_INV
    );
  TD1_TRIAC_TRIG_I_D2_PT_3_0_INV_763 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => TD1_TRIAC_TRIG_I_D2_PT_3_0_INV
    );
  TD1_TRIAC_TRIG_I_D2_PT_4_0_INV_764 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => TD1_TRIAC_TRIG_I_D2_PT_4_0_INV
    );
  TD1_TRIAC_TRIG_I_XOR_0_INV_765 : X_INV 
    port map (
      I => TD1_TRIAC_TRIG_I_D1,
      O => TD1_TRIAC_TRIG_I_XOR_0_INV
    );
  EXP1_EXP_PT_0_0_INV_766 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => EXP1_EXP_PT_0_0_INV
    );
  EXP1_EXP_PT_0_1_INV_767 : X_INV 
    port map (
      I => LIGHT_VALUE(5),
      O => EXP1_EXP_PT_0_1_INV
    );
  EXP1_EXP_PT_1_0_INV_768 : X_INV 
    port map (
      I => LIGHT_VALUE(5),
      O => EXP1_EXP_PT_1_0_INV
    );
  LIGHT_VALUE_4_RSTF_PT_0_0_INV_769 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => LIGHT_VALUE_4_RSTF_PT_0_0_INV
    );
  LIGHT_VALUE_4_RSTF_PT_0_1_INV_770 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => LIGHT_VALUE_4_RSTF_PT_0_1_INV
    );
  LIGHT_VALUE_4_D2_PT_1_8_INV_771 : X_INV 
    port map (
      I => LIGHT_VALUE(5),
      O => LIGHT_VALUE_4_D2_PT_1_8_INV
    );
  LIGHT_VALUE_4_D2_PT_1_12_INV_772 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => LIGHT_VALUE_4_D2_PT_1_12_INV
    );
  LIGHT_VALUE_4_EXP_PT_0_0_INV_773 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => LIGHT_VALUE_4_EXP_PT_0_0_INV
    );
  LIGHT_VALUE_4_EXP_PT_0_2_INV_774 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => LIGHT_VALUE_4_EXP_PT_0_2_INV
    );
  LIGHT_VALUE_4_EXP_PT_0_3_INV_775 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => LIGHT_VALUE_4_EXP_PT_0_3_INV
    );
  LIGHT_VALUE_4_EXP_PT_0_4_INV_776 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => LIGHT_VALUE_4_EXP_PT_0_4_INV
    );
  LIGHT_VALUE_4_EXP_PT_0_5_INV_777 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => LIGHT_VALUE_4_EXP_PT_0_5_INV
    );
  LIGHT_VALUE_4_EXP_PT_1_0_INV_778 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => LIGHT_VALUE_4_EXP_PT_1_0_INV
    );
  LIGHT_VALUE_4_EXP_PT_1_1_INV_779 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => LIGHT_VALUE_4_EXP_PT_1_1_INV
    );
  LIGHT_VALUE_4_EXP_PT_1_2_INV_780 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => LIGHT_VALUE_4_EXP_PT_1_2_INV
    );
  LIGHT_VALUE_4_EXP_PT_1_3_INV_781 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => LIGHT_VALUE_4_EXP_PT_1_3_INV
    );
  LIGHT_VALUE_4_EXP_PT_1_4_INV_782 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => LIGHT_VALUE_4_EXP_PT_1_4_INV
    );
  LIGHT_VALUE_4_EXP_PT_2_1_INV_783 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => LIGHT_VALUE_4_EXP_PT_2_1_INV
    );
  LIGHT_VALUE_4_EXP_PT_2_6_INV_784 : X_INV 
    port map (
      I => LIGHT_VALUE(3),
      O => LIGHT_VALUE_4_EXP_PT_2_6_INV
    );
  LIGHT_VALUE_4_EXP_PT_2_7_INV_785 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => LIGHT_VALUE_4_EXP_PT_2_7_INV
    );
  EXP0_EXP_PT_0_0_INV_786 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP0_EXP_PT_0_0_INV
    );
  EXP0_EXP_PT_0_2_INV_787 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP0_EXP_PT_0_2_INV
    );
  EXP0_EXP_PT_0_3_INV_788 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP0_EXP_PT_0_3_INV
    );
  EXP0_EXP_PT_0_4_INV_789 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP0_EXP_PT_0_4_INV
    );
  EXP0_EXP_PT_0_5_INV_790 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP0_EXP_PT_0_5_INV
    );
  EXP0_EXP_PT_0_6_INV_791 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => EXP0_EXP_PT_0_6_INV
    );
  EXP0_EXP_PT_0_7_INV_792 : X_INV 
    port map (
      I => FC1_CNT_6_FBK,
      O => EXP0_EXP_PT_0_7_INV
    );
  EXP0_EXP_PT_0_8_INV_793 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP0_EXP_PT_0_8_INV
    );
  EXP0_EXP_PT_0_9_INV_794 : X_INV 
    port map (
      I => LIGHT_VALUE(3),
      O => EXP0_EXP_PT_0_9_INV
    );
  EXP0_EXP_PT_0_10_INV_795 : X_INV 
    port map (
      I => LIGHT_VALUE(1),
      O => EXP0_EXP_PT_0_10_INV
    );
  EXP0_EXP_PT_0_11_INV_796 : X_INV 
    port map (
      I => LIGHT_VALUE(2),
      O => EXP0_EXP_PT_0_11_INV
    );
  EXP0_EXP_PT_0_13_INV_797 : X_INV 
    port map (
      I => LIGHT_VALUE(0),
      O => EXP0_EXP_PT_0_13_INV
    );
  EXP0_EXP_PT_0_14_INV_798 : X_INV 
    port map (
      I => FC1_CNT_7_FBK,
      O => EXP0_EXP_PT_0_14_INV
    );
  EXP0_EXP_PT_1_0_INV_799 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP0_EXP_PT_1_0_INV
    );
  EXP0_EXP_PT_1_1_INV_800 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP0_EXP_PT_1_1_INV
    );
  EXP0_EXP_PT_1_2_INV_801 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP0_EXP_PT_1_2_INV
    );
  EXP0_EXP_PT_1_3_INV_802 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP0_EXP_PT_1_3_INV
    );
  EXP0_EXP_PT_1_4_INV_803 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP0_EXP_PT_1_4_INV
    );
  EXP0_EXP_PT_1_5_INV_804 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => EXP0_EXP_PT_1_5_INV
    );
  EXP0_EXP_PT_1_6_INV_805 : X_INV 
    port map (
      I => FC1_CNT_6_FBK,
      O => EXP0_EXP_PT_1_6_INV
    );
  EXP0_EXP_PT_1_7_INV_806 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP0_EXP_PT_1_7_INV
    );
  EXP0_EXP_PT_1_9_INV_807 : X_INV 
    port map (
      I => LIGHT_VALUE(3),
      O => EXP0_EXP_PT_1_9_INV
    );
  EXP0_EXP_PT_1_10_INV_808 : X_INV 
    port map (
      I => LIGHT_VALUE(1),
      O => EXP0_EXP_PT_1_10_INV
    );
  EXP0_EXP_PT_1_11_INV_809 : X_INV 
    port map (
      I => LIGHT_VALUE(2),
      O => EXP0_EXP_PT_1_11_INV
    );
  EXP0_EXP_PT_1_13_INV_810 : X_INV 
    port map (
      I => LIGHT_VALUE(0),
      O => EXP0_EXP_PT_1_13_INV
    );
  EXP0_EXP_PT_1_14_INV_811 : X_INV 
    port map (
      I => FC1_CNT_7_FBK,
      O => EXP0_EXP_PT_1_14_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_0_1_INV_812 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_0_1_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_1_1_INV_813 : X_INV 
    port map (
      I => CM_PANIC_ON,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_1_1_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_1_2_INV_814 : X_INV 
    port map (
      I => CM_FADE_UP,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_1_2_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_1_INV_815 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_1_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_5_INV_816 : X_INV 
    port map (
      I => LIGHT_VALUE(2),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_5_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_6_INV_817 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_6_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_7_INV_818 : X_INV 
    port map (
      I => LIGHT_VALUE(0),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_2_7_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_0_INV_819 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_0_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_1_INV_820 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_1_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_2_INV_821 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_2_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_3_INV_822 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_3_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_4_INV_823 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_4_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_5_INV_824 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_5_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_6_INV_825 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_6_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_7_INV_826 : X_INV 
    port map (
      I => FC1_CNT_6_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_7_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_8_INV_827 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_8_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_9_INV_828 : X_INV 
    port map (
      I => LIGHT_VALUE(5),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_9_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_10_INV_829 : X_INV 
    port map (
      I => LIGHT_VALUE(3),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_10_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_11_INV_830 : X_INV 
    port map (
      I => LIGHT_VALUE(1),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_11_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_12_INV_831 : X_INV 
    port map (
      I => LIGHT_VALUE(2),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_12_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_14_INV_832 : X_INV 
    port map (
      I => CM_PANIC_ON,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_14_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_15_INV_833 : X_INV 
    port map (
      I => LIGHT_VALUE(0),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_15_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_16_INV_834 : X_INV 
    port map (
      I => FC1_CNT_7_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_EXP_PT_3_16_INV
    );
  EXP2_EXP_PT_0_2_INV_835 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP2_EXP_PT_0_2_INV
    );
  EXP2_EXP_PT_1_0_INV_836 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP2_EXP_PT_1_0_INV
    );
  EXP2_EXP_PT_1_2_INV_837 : X_INV 
    port map (
      I => CM_PANIC_ON,
      O => EXP2_EXP_PT_1_2_INV
    );
  EXP2_EXP_PT_2_1_INV_838 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => EXP2_EXP_PT_2_1_INV
    );
  EXP2_EXP_PT_2_5_INV_839 : X_INV 
    port map (
      I => LIGHT_VALUE(2),
      O => EXP2_EXP_PT_2_5_INV
    );
  EXP2_EXP_PT_2_6_INV_840 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP2_EXP_PT_2_6_INV
    );
  EXP2_EXP_PT_2_7_INV_841 : X_INV 
    port map (
      I => LIGHT_VALUE(0),
      O => EXP2_EXP_PT_2_7_INV
    );
  EXP2_EXP_PT_3_0_INV_842 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP2_EXP_PT_3_0_INV
    );
  EXP2_EXP_PT_3_1_INV_843 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => EXP2_EXP_PT_3_1_INV
    );
  EXP2_EXP_PT_3_2_INV_844 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP2_EXP_PT_3_2_INV
    );
  EXP2_EXP_PT_3_3_INV_845 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP2_EXP_PT_3_3_INV
    );
  EXP2_EXP_PT_3_4_INV_846 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP2_EXP_PT_3_4_INV
    );
  EXP2_EXP_PT_3_5_INV_847 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP2_EXP_PT_3_5_INV
    );
  EXP2_EXP_PT_3_6_INV_848 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => EXP2_EXP_PT_3_6_INV
    );
  EXP2_EXP_PT_3_7_INV_849 : X_INV 
    port map (
      I => FC1_CNT_6_FBK,
      O => EXP2_EXP_PT_3_7_INV
    );
  EXP2_EXP_PT_3_8_INV_850 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP2_EXP_PT_3_8_INV
    );
  EXP2_EXP_PT_3_9_INV_851 : X_INV 
    port map (
      I => LIGHT_VALUE(5),
      O => EXP2_EXP_PT_3_9_INV
    );
  EXP2_EXP_PT_3_10_INV_852 : X_INV 
    port map (
      I => LIGHT_VALUE(3),
      O => EXP2_EXP_PT_3_10_INV
    );
  EXP2_EXP_PT_3_11_INV_853 : X_INV 
    port map (
      I => LIGHT_VALUE(1),
      O => EXP2_EXP_PT_3_11_INV
    );
  EXP2_EXP_PT_3_12_INV_854 : X_INV 
    port map (
      I => LIGHT_VALUE(2),
      O => EXP2_EXP_PT_3_12_INV
    );
  EXP2_EXP_PT_3_14_INV_855 : X_INV 
    port map (
      I => CM_PANIC_ON,
      O => EXP2_EXP_PT_3_14_INV
    );
  EXP2_EXP_PT_3_15_INV_856 : X_INV 
    port map (
      I => LIGHT_VALUE(0),
      O => EXP2_EXP_PT_3_15_INV
    );
  EXP2_EXP_PT_3_16_INV_857 : X_INV 
    port map (
      I => FC1_CNT_7_FBK,
      O => EXP2_EXP_PT_3_16_INV
    );
  CM_FADE_DOWN_D2_PT_2_0_INV_858 : X_INV 
    port map (
      I => RXD_READY_FBK,
      O => CM_FADE_DOWN_D2_PT_2_0_INV
    );
  CM_FADE_DOWN_D2_PT_2_1_INV_859 : X_INV 
    port map (
      I => RXD_READY_FBK,
      O => CM_FADE_DOWN_D2_PT_2_1_INV
    );
  CM_FADE_DOWN_D2_PT_5_1_INV_860 : X_INV 
    port map (
      I => RXD_4_FBK,
      O => CM_FADE_DOWN_D2_PT_5_1_INV
    );
  CM_FADE_DOWN_D2_PT_6_0_INV_861 : X_INV 
    port map (
      I => RC_ADDRESS_C(0),
      O => CM_FADE_DOWN_D2_PT_6_0_INV
    );
  CM_FADE_DOWN_XOR_0_INV_862 : X_INV 
    port map (
      I => CM_FADE_DOWN_D1,
      O => CM_FADE_DOWN_XOR_0_INV
    );
  RXD_READY_EXP_PT_0_1_INV_863 : X_INV 
    port map (
      I => RXD_5_FBK,
      O => RXD_READY_EXP_PT_0_1_INV
    );
  RXD_READY_EXP_PT_1_0_INV_864 : X_INV 
    port map (
      I => RC_ADDRESS_C(1),
      O => RXD_READY_EXP_PT_1_0_INV
    );
  RXD_READY_EXP_PT_2_1_INV_865 : X_INV 
    port map (
      I => RXD_6_FBK,
      O => RXD_READY_EXP_PT_2_1_INV
    );
  RXD_READY_EXP_PT_3_0_INV_866 : X_INV 
    port map (
      I => RC_ADDRESS_C(2),
      O => RXD_READY_EXP_PT_3_0_INV
    );
  RXD_READY_EXP_PT_4_1_INV_867 : X_INV 
    port map (
      I => RXD_7_FBK,
      O => RXD_READY_EXP_PT_4_1_INV
    );
  RXD_7_EXP_PT_0_1_INV_868 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_7_EXP_PT_0_1_INV
    );
  RXD_7_EXP_PT_1_0_INV_869 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_7_EXP_PT_1_0_INV
    );
  RXD_7_D2_PT_0_1_INV_870 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_7_D2_PT_0_1_INV
    );
  RXD_7_D2_PT_0_3_INV_871 : X_INV 
    port map (
      I => UAR1_BYTE_OUT(7),
      O => RXD_7_D2_PT_0_3_INV
    );
  RXD_7_D2_PT_1_1_INV_872 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_7_D2_PT_1_1_INV
    );
  RXD_7_D2_PT_1_2_INV_873 : X_INV 
    port map (
      I => RXD_7_FBK,
      O => RXD_7_D2_PT_1_2_INV
    );
  UAR1_BYTE_AVAIL_D2_PT_0_2_INV_874 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS_0_FBK,
      O => UAR1_BYTE_AVAIL_D2_PT_0_2_INV
    );
  UAR1_BYTE_AVAIL_D2_PT_0_3_INV_875 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS_1_FBK,
      O => UAR1_BYTE_AVAIL_D2_PT_0_3_INV
    );
  UAR1_BYTE_AVAIL_D2_PT_0_4_INV_876 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS_2_FBK,
      O => UAR1_BYTE_AVAIL_D2_PT_0_4_INV
    );
  UAR1_BIT_DONE_D2_PT_0_0_INV_877 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL_FBK,
      O => UAR1_BIT_DONE_D2_PT_0_0_INV
    );
  UAR1_BIT_DONE_D2_PT_0_1_INV_878 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_Q_5,
      O => UAR1_BIT_DONE_D2_PT_0_1_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_2_0_INV_879 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_2_0_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_2_2_INV_880 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_2_2_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_2_3_INV_881 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_2_3_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_2_4_INV_882 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_2_4_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_2_5_INV_883 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q_6,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_2_5_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_2_6_INV_884 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_FBK,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_2_6_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_3_0_INV_885 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_3_0_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_3_1_INV_886 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_3_1_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_3_2_INV_887 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_3_2_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_3_3_INV_888 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_3_3_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_3_5_INV_889 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q_6,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_3_5_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_3_6_INV_890 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_FBK,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_3_6_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_4_0_INV_891 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_4_0_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_4_1_INV_892 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_4_1_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_4_2_INV_893 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_4_2_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_4_3_INV_894 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_4_3_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_4_5_INV_895 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q_6,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_4_5_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_4_6_INV_896 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_FBK,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_4_6_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_5_0_INV_897 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_5_0_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_5_1_INV_898 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_5_1_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_5_2_INV_899 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_5_2_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_5_3_INV_900 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_5_3_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_5_5_INV_901 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q_6,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_5_5_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_5_6_INV_902 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_FBK,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_5_6_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_6_0_INV_903 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_6_0_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_6_1_INV_904 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_6_1_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_6_2_INV_905 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_6_2_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_6_3_INV_906 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_6_3_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_6_5_INV_907 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q_6,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_6_5_INV
    );
  UAR1_BC1_CURRENT_STATE_11_D2_PT_6_6_INV_908 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_FBK,
      O => UAR1_BC1_CURRENT_STATE_11_D2_PT_6_6_INV
    );
  UAR1_BC1_CURRENT_STATE_11_XOR_0_INV_909 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_D1,
      O => UAR1_BC1_CURRENT_STATE_11_XOR_0_INV
    );
  EXP9_EXP_PT_0_1_INV_910 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => EXP9_EXP_PT_0_1_INV
    );
  EXP9_EXP_PT_0_5_INV_911 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_1_FBK,
      O => EXP9_EXP_PT_0_5_INV
    );
  EXP9_EXP_PT_1_1_INV_912 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => EXP9_EXP_PT_1_1_INV
    );
  EXP9_EXP_PT_1_2_INV_913 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => EXP9_EXP_PT_1_2_INV
    );
  EXP9_EXP_PT_1_3_INV_914 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => EXP9_EXP_PT_1_3_INV
    );
  EXP9_EXP_PT_1_4_INV_915 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => EXP9_EXP_PT_1_4_INV
    );
  EXP9_EXP_PT_1_5_INV_916 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q_6,
      O => EXP9_EXP_PT_1_5_INV
    );
  EXP9_EXP_PT_2_0_INV_917 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => EXP9_EXP_PT_2_0_INV
    );
  EXP9_EXP_PT_2_4_INV_918 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_1_FBK,
      O => EXP9_EXP_PT_2_4_INV
    );
  EXP9_EXP_PT_2_5_INV_919 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_FBK,
      O => EXP9_EXP_PT_2_5_INV
    );
  EXP9_EXP_PT_3_0_INV_920 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => EXP9_EXP_PT_3_0_INV
    );
  EXP9_EXP_PT_3_1_INV_921 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => EXP9_EXP_PT_3_1_INV
    );
  EXP9_EXP_PT_3_2_INV_922 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => EXP9_EXP_PT_3_2_INV
    );
  EXP9_EXP_PT_3_3_INV_923 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => EXP9_EXP_PT_3_3_INV
    );
  EXP9_EXP_PT_3_4_INV_924 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q_6,
      O => EXP9_EXP_PT_3_4_INV
    );
  EXP9_EXP_PT_3_6_INV_925 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_FBK,
      O => EXP9_EXP_PT_3_6_INV
    );
  EXP9_EXP_PT_4_1_INV_926 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => EXP9_EXP_PT_4_1_INV
    );
  EXP9_EXP_PT_4_2_INV_927 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_3_FBK,
      O => EXP9_EXP_PT_4_2_INV
    );
  EXP9_EXP_PT_4_3_INV_928 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_2_FBK,
      O => EXP9_EXP_PT_4_3_INV
    );
  EXP9_EXP_PT_4_4_INV_929 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_4_FBK,
      O => EXP9_EXP_PT_4_4_INV
    );
  EXP9_EXP_PT_4_5_INV_930 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_5_FBK,
      O => EXP9_EXP_PT_4_5_INV
    );
  EXP9_EXP_PT_4_6_INV_931 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_6_FBK,
      O => EXP9_EXP_PT_4_6_INV
    );
  EXP9_EXP_PT_4_7_INV_932 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_7_FBK,
      O => EXP9_EXP_PT_4_7_INV
    );
  EXP9_EXP_PT_4_8_INV_933 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_8_FBK,
      O => EXP9_EXP_PT_4_8_INV
    );
  EXP9_EXP_PT_4_9_INV_934 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_9_FBK,
      O => EXP9_EXP_PT_4_9_INV
    );
  EXP9_EXP_PT_4_10_INV_935 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q_6,
      O => EXP9_EXP_PT_4_10_INV
    );
  EXP9_EXP_PT_4_11_INV_936 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_1_FBK,
      O => EXP9_EXP_PT_4_11_INV
    );
  UAR1_BM1_SAMPLED_BITS_0_D2_PT_1_0_INV_937 : X_INV 
    port map (
      I => UAR1_BM1_CURRENT_STATE_3_FBK,
      O => UAR1_BM1_SAMPLED_BITS_0_D2_PT_1_0_INV
    );
  UAR1_BM1_CURRENT_STATE_3_D2_PT_0_0_INV_938 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL_FBK,
      O => UAR1_BM1_CURRENT_STATE_3_D2_PT_0_0_INV
    );
  UAR1_BM1_CURRENT_STATE_3_D2_PT_0_1_INV_939 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_Q_5,
      O => UAR1_BM1_CURRENT_STATE_3_D2_PT_0_1_INV
    );
  UAR1_BM1_CURRENT_STATE_3_D2_PT_1_0_INV_940 : X_INV 
    port map (
      I => UAR1_BIT_DONE_FBK,
      O => UAR1_BM1_CURRENT_STATE_3_D2_PT_1_0_INV
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_0_0_INV_941 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL_FBK,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_0_0_INV
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_0_1_INV_942 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_Q_5,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_0_1_INV
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_0_INV_943 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL_FBK,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_0_INV
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_1_INV_944 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_Q_5,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_1_INV
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_2_INV_945 : X_INV 
    port map (
      I => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_FBK,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_1_2_INV
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_0_INV_946 : X_INV 
    port map (
      I => UAR1_BM1_CURRENT_STATE_1_FBK,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_0_INV
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_1_INV_947 : X_INV 
    port map (
      I => UAR1_BIT_DONE_FBK,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_1_INV
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_3_INV_948 : X_INV 
    port map (
      I => UAR1_BM1_CURRENT_STATE_2_FBK,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_3_INV
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_4_INV_949 : X_INV 
    port map (
      I => UAR1_BM1_CURRENT_STATE_3_FBK,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D2_PT_2_4_INV
    );
  UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_XOR_0_INV_950 : X_INV 
    port map (
      I => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_D1,
      O => UAR1_BM1_CURRENT_STATE_H_CURRENT_STATE_4_XOR_0_INV
    );
  UAR1_BM1_CURRENT_STATE_1_D2_PT_0_0_INV_951 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL_FBK,
      O => UAR1_BM1_CURRENT_STATE_1_D2_PT_0_0_INV
    );
  UAR1_BM1_CURRENT_STATE_1_D2_PT_0_1_INV_952 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_Q_5,
      O => UAR1_BM1_CURRENT_STATE_1_D2_PT_0_1_INV
    );
  UAR1_BM1_CURRENT_STATE_2_D2_PT_0_0_INV_953 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL_FBK,
      O => UAR1_BM1_CURRENT_STATE_2_D2_PT_0_0_INV
    );
  UAR1_BM1_CURRENT_STATE_2_D2_PT_0_1_INV_954 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_Q_5,
      O => UAR1_BM1_CURRENT_STATE_2_D2_PT_0_1_INV
    );
  UAR1_BM1_SAMPLED_BITS_1_D2_PT_1_0_INV_955 : X_INV 
    port map (
      I => UAR1_BM1_CURRENT_STATE_2_FBK,
      O => UAR1_BM1_SAMPLED_BITS_1_D2_PT_1_0_INV
    );
  UAR1_BM1_SAMPLED_BITS_2_D2_PT_1_0_INV_956 : X_INV 
    port map (
      I => UAR1_BM1_CURRENT_STATE_1_FBK,
      O => UAR1_BM1_SAMPLED_BITS_2_D2_PT_1_0_INV
    );
  UAR1_BC1_CURRENT_STATE_1_D2_PT_0_0_INV_957 : X_INV 
    port map (
      I => UAR1_BIT_DONE,
      O => UAR1_BC1_CURRENT_STATE_1_D2_PT_0_0_INV
    );
  UAR1_BC1_CURRENT_STATE_1_D2_PT_2_1_INV_958 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_1_D2_PT_2_1_INV
    );
  UAR1_BC1_CURRENT_STATE_1_D2_PT_2_2_INV_959 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_1_D2_PT_2_2_INV
    );
  UAR1_BC1_CURRENT_STATE_1_D2_PT_2_3_INV_960 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_1_D2_PT_2_3_INV
    );
  UAR1_BC1_CURRENT_STATE_2_D2_PT_0_0_INV_961 : X_INV 
    port map (
      I => UAR1_BIT_DONE,
      O => UAR1_BC1_CURRENT_STATE_2_D2_PT_0_0_INV
    );
  UAR1_BC1_CURRENT_STATE_2_D2_PT_2_2_INV_962 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_2_D2_PT_2_2_INV
    );
  UAR1_BC1_CURRENT_STATE_2_D2_PT_2_3_INV_963 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_2_D2_PT_2_3_INV
    );
  UAR1_BC1_CURRENT_STATE_2_D2_PT_2_4_INV_964 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_2_D2_PT_2_4_INV
    );
  UAR1_BC1_CURRENT_STATE_3_D2_PT_0_0_INV_965 : X_INV 
    port map (
      I => UAR1_BIT_DONE,
      O => UAR1_BC1_CURRENT_STATE_3_D2_PT_0_0_INV
    );
  UAR1_BC1_CURRENT_STATE_3_D2_PT_2_1_INV_966 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_3_D2_PT_2_1_INV
    );
  UAR1_BC1_CURRENT_STATE_3_D2_PT_2_2_INV_967 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_3_D2_PT_2_2_INV
    );
  UAR1_BC1_CURRENT_STATE_3_D2_PT_2_3_INV_968 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_3_D2_PT_2_3_INV
    );
  UAR1_BC1_CURRENT_STATE_4_D2_PT_0_0_INV_969 : X_INV 
    port map (
      I => UAR1_BIT_DONE,
      O => UAR1_BC1_CURRENT_STATE_4_D2_PT_0_0_INV
    );
  UAR1_BC1_CURRENT_STATE_4_D2_PT_2_1_INV_970 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_4_D2_PT_2_1_INV
    );
  UAR1_BC1_CURRENT_STATE_4_D2_PT_2_2_INV_971 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_4_D2_PT_2_2_INV
    );
  UAR1_BC1_CURRENT_STATE_4_D2_PT_2_3_INV_972 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_4_D2_PT_2_3_INV
    );
  UAR1_BC1_CURRENT_STATE_5_D2_PT_0_0_INV_973 : X_INV 
    port map (
      I => UAR1_BIT_DONE,
      O => UAR1_BC1_CURRENT_STATE_5_D2_PT_0_0_INV
    );
  UAR1_BC1_CURRENT_STATE_5_D2_PT_2_1_INV_974 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_5_D2_PT_2_1_INV
    );
  UAR1_BC1_CURRENT_STATE_5_D2_PT_2_2_INV_975 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_5_D2_PT_2_2_INV
    );
  UAR1_BC1_CURRENT_STATE_5_D2_PT_2_3_INV_976 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_5_D2_PT_2_3_INV
    );
  UAR1_BC1_CURRENT_STATE_6_D2_PT_0_0_INV_977 : X_INV 
    port map (
      I => UAR1_BIT_DONE,
      O => UAR1_BC1_CURRENT_STATE_6_D2_PT_0_0_INV
    );
  UAR1_BC1_CURRENT_STATE_6_D2_PT_2_1_INV_978 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_6_D2_PT_2_1_INV
    );
  UAR1_BC1_CURRENT_STATE_6_D2_PT_2_2_INV_979 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_6_D2_PT_2_2_INV
    );
  UAR1_BC1_CURRENT_STATE_6_D2_PT_2_3_INV_980 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_6_D2_PT_2_3_INV
    );
  UAR1_BC1_CURRENT_STATE_7_D2_PT_0_0_INV_981 : X_INV 
    port map (
      I => UAR1_BIT_DONE,
      O => UAR1_BC1_CURRENT_STATE_7_D2_PT_0_0_INV
    );
  UAR1_BC1_CURRENT_STATE_7_D2_PT_2_1_INV_982 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_7_D2_PT_2_1_INV
    );
  UAR1_BC1_CURRENT_STATE_7_D2_PT_2_2_INV_983 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_7_D2_PT_2_2_INV
    );
  UAR1_BC1_CURRENT_STATE_7_D2_PT_2_3_INV_984 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_7_D2_PT_2_3_INV
    );
  UAR1_BC1_CURRENT_STATE_8_D2_PT_0_0_INV_985 : X_INV 
    port map (
      I => UAR1_BIT_DONE,
      O => UAR1_BC1_CURRENT_STATE_8_D2_PT_0_0_INV
    );
  UAR1_BC1_CURRENT_STATE_8_D2_PT_2_1_INV_986 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => UAR1_BC1_CURRENT_STATE_8_D2_PT_2_1_INV
    );
  UAR1_BC1_CURRENT_STATE_8_D2_PT_2_2_INV_987 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => UAR1_BC1_CURRENT_STATE_8_D2_PT_2_2_INV
    );
  UAR1_BC1_CURRENT_STATE_8_D2_PT_2_3_INV_988 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => UAR1_BC1_CURRENT_STATE_8_D2_PT_2_3_INV
    );
  UAR1_BC1_CURRENT_STATE_9_D2_PT_0_0_INV_989 : X_INV 
    port map (
      I => UAR1_BIT_DONE,
      O => UAR1_BC1_CURRENT_STATE_9_D2_PT_0_0_INV
    );
  UAR1_BC1_CURRENT_STATE_10_D2_PT_1_0_INV_990 : X_INV 
    port map (
      I => UAR1_BIT_DONE_FBK,
      O => UAR1_BC1_CURRENT_STATE_10_D2_PT_1_0_INV
    );
  EXP10_EXP_PT_0_0_INV_991 : X_INV 
    port map (
      I => UAR1_BIT_DONE,
      O => EXP10_EXP_PT_0_0_INV
    );
  EXP10_EXP_PT_0_2_INV_992 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => EXP10_EXP_PT_0_2_INV
    );
  EXP10_EXP_PT_1_0_INV_993 : X_INV 
    port map (
      I => UAR1_BIT_DONE,
      O => EXP10_EXP_PT_1_0_INV
    );
  EXP10_EXP_PT_1_1_INV_994 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => EXP10_EXP_PT_1_1_INV
    );
  EXP10_EXP_PT_1_2_INV_995 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_FBK,
      O => EXP10_EXP_PT_1_2_INV
    );
  EXP10_EXP_PT_2_0_INV_996 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => EXP10_EXP_PT_2_0_INV
    );
  EXP10_EXP_PT_2_1_INV_997 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => EXP10_EXP_PT_2_1_INV
    );
  EXP10_EXP_PT_2_2_INV_998 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => EXP10_EXP_PT_2_2_INV
    );
  EXP10_EXP_PT_2_3_INV_999 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => EXP10_EXP_PT_2_3_INV
    );
  EXP10_EXP_PT_2_5_INV_1000 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q_6,
      O => EXP10_EXP_PT_2_5_INV
    );
  EXP10_EXP_PT_2_6_INV_1001 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_FBK,
      O => EXP10_EXP_PT_2_6_INV
    );
  EXP10_EXP_PT_3_0_INV_1002 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => EXP10_EXP_PT_3_0_INV
    );
  EXP10_EXP_PT_3_1_INV_1003 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => EXP10_EXP_PT_3_1_INV
    );
  EXP10_EXP_PT_3_2_INV_1004 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => EXP10_EXP_PT_3_2_INV
    );
  EXP10_EXP_PT_3_3_INV_1005 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => EXP10_EXP_PT_3_3_INV
    );
  EXP10_EXP_PT_3_5_INV_1006 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q_6,
      O => EXP10_EXP_PT_3_5_INV
    );
  EXP10_EXP_PT_3_6_INV_1007 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_FBK,
      O => EXP10_EXP_PT_3_6_INV
    );
  EXP10_EXP_PT_4_0_INV_1008 : X_INV 
    port map (
      I => UAR1_BYTE_AVAIL,
      O => EXP10_EXP_PT_4_0_INV
    );
  EXP10_EXP_PT_4_1_INV_1009 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(0),
      O => EXP10_EXP_PT_4_1_INV
    );
  EXP10_EXP_PT_4_2_INV_1010 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(1),
      O => EXP10_EXP_PT_4_2_INV
    );
  EXP10_EXP_PT_4_3_INV_1011 : X_INV 
    port map (
      I => UAR1_BM1_SAMPLED_BITS(2),
      O => EXP10_EXP_PT_4_3_INV
    );
  EXP10_EXP_PT_4_5_INV_1012 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_10_Q_6,
      O => EXP10_EXP_PT_4_5_INV
    );
  EXP10_EXP_PT_4_6_INV_1013 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_11_FBK,
      O => EXP10_EXP_PT_4_6_INV
    );
  UAR1_BYTE_OUT_7_D2_PT_0_0_INV_1014 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_2_Q_7,
      O => UAR1_BYTE_OUT_7_D2_PT_0_0_INV
    );
  RXD_5_D2_PT_0_1_INV_1015 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_5_D2_PT_0_1_INV
    );
  RXD_5_D2_PT_0_3_INV_1016 : X_INV 
    port map (
      I => UAR1_BYTE_OUT(5),
      O => RXD_5_D2_PT_0_3_INV
    );
  RXD_5_D2_PT_1_1_INV_1017 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_5_D2_PT_1_1_INV
    );
  RXD_5_D2_PT_1_2_INV_1018 : X_INV 
    port map (
      I => RXD_5_FBK,
      O => RXD_5_D2_PT_1_2_INV
    );
  UAR1_BYTE_OUT_5_D2_PT_0_0_INV_1019 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_4_FBK,
      O => UAR1_BYTE_OUT_5_D2_PT_0_0_INV
    );
  RXD_6_D2_PT_0_1_INV_1020 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_6_D2_PT_0_1_INV
    );
  RXD_6_D2_PT_0_3_INV_1021 : X_INV 
    port map (
      I => UAR1_BYTE_OUT(6),
      O => RXD_6_D2_PT_0_3_INV
    );
  RXD_6_D2_PT_1_1_INV_1022 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_6_D2_PT_1_1_INV
    );
  RXD_6_D2_PT_1_2_INV_1023 : X_INV 
    port map (
      I => RXD_6_FBK,
      O => RXD_6_D2_PT_1_2_INV
    );
  UAR1_BYTE_OUT_6_D2_PT_0_0_INV_1024 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_3_Q_8,
      O => UAR1_BYTE_OUT_6_D2_PT_0_0_INV
    );
  RXD_2_D2_PT_0_1_INV_1025 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_2_D2_PT_0_1_INV
    );
  RXD_2_D2_PT_0_3_INV_1026 : X_INV 
    port map (
      I => UAR1_BYTE_OUT(2),
      O => RXD_2_D2_PT_0_3_INV
    );
  RXD_2_D2_PT_1_1_INV_1027 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_2_D2_PT_1_1_INV
    );
  RXD_2_D2_PT_1_2_INV_1028 : X_INV 
    port map (
      I => RXD_2_FBK,
      O => RXD_2_D2_PT_1_2_INV
    );
  UAR1_BYTE_OUT_2_D2_PT_0_0_INV_1029 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_7_FBK,
      O => UAR1_BYTE_OUT_2_D2_PT_0_0_INV
    );
  EXP19_EXP_PT_0_1_INV_1030 : X_INV 
    port map (
      I => RXD_5_FBK,
      O => EXP19_EXP_PT_0_1_INV
    );
  EXP19_EXP_PT_1_0_INV_1031 : X_INV 
    port map (
      I => RC_ADDRESS_C(1),
      O => EXP19_EXP_PT_1_0_INV
    );
  EXP19_EXP_PT_2_1_INV_1032 : X_INV 
    port map (
      I => RXD_6_FBK,
      O => EXP19_EXP_PT_2_1_INV
    );
  EXP19_EXP_PT_3_0_INV_1033 : X_INV 
    port map (
      I => RC_ADDRESS_C(2),
      O => EXP19_EXP_PT_3_0_INV
    );
  EXP19_EXP_PT_4_1_INV_1034 : X_INV 
    port map (
      I => RXD_7_FBK,
      O => EXP19_EXP_PT_4_1_INV
    );
  EXP20_EXP_PT_1_1_INV_1035 : X_INV 
    port map (
      I => CM_FADE_DOWN_FBK,
      O => EXP20_EXP_PT_1_1_INV
    );
  EXP20_EXP_PT_3_0_INV_1036 : X_INV 
    port map (
      I => CM_FADE_DOWN_FBK,
      O => EXP20_EXP_PT_3_0_INV
    );
  EXP20_EXP_PT_4_0_INV_1037 : X_INV 
    port map (
      I => CM_FADE_DOWN_FBK,
      O => EXP20_EXP_PT_4_0_INV
    );
  EXP20_EXP_PT_4_1_INV_1038 : X_INV 
    port map (
      I => RXD_0_FBK,
      O => EXP20_EXP_PT_4_1_INV
    );
  EXP20_EXP_PT_5_0_INV_1039 : X_INV 
    port map (
      I => RC_ADDRESS_C(3),
      O => EXP20_EXP_PT_5_0_INV
    );
  RXD_1_EXP_PT_1_0_INV_1040 : X_INV 
    port map (
      I => RXD_3_FBK,
      O => RXD_1_EXP_PT_1_0_INV
    );
  RXD_1_EXP_PT_1_2_INV_1041 : X_INV 
    port map (
      I => RXD_1_FBK,
      O => RXD_1_EXP_PT_1_2_INV
    );
  RXD_1_D2_PT_0_1_INV_1042 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_1_D2_PT_0_1_INV
    );
  RXD_1_D2_PT_0_3_INV_1043 : X_INV 
    port map (
      I => RXD_1_FBK,
      O => RXD_1_D2_PT_0_3_INV
    );
  RXD_1_D2_PT_1_1_INV_1044 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_1_D2_PT_1_1_INV
    );
  RXD_1_D2_PT_1_2_INV_1045 : X_INV 
    port map (
      I => UAR1_BYTE_OUT(1),
      O => RXD_1_D2_PT_1_2_INV
    );
  UAR1_BYTE_OUT_1_D2_PT_0_0_INV_1046 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_8_FBK,
      O => UAR1_BYTE_OUT_1_D2_PT_0_0_INV
    );
  RXD_3_D2_PT_0_2_INV_1047 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_3_D2_PT_0_2_INV
    );
  RXD_3_D2_PT_0_3_INV_1048 : X_INV 
    port map (
      I => UAR1_BYTE_OUT(3),
      O => RXD_3_D2_PT_0_3_INV
    );
  RXD_3_D2_PT_1_0_INV_1049 : X_INV 
    port map (
      I => RXD_3_FBK,
      O => RXD_3_D2_PT_1_0_INV
    );
  RXD_3_D2_PT_1_2_INV_1050 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_3_D2_PT_1_2_INV
    );
  UAR1_BYTE_OUT_3_D2_PT_0_0_INV_1051 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_6_FBK,
      O => UAR1_BYTE_OUT_3_D2_PT_0_0_INV
    );
  RXD_0_EXP_PT_1_0_INV_1052 : X_INV 
    port map (
      I => RXD_1_FBK,
      O => RXD_0_EXP_PT_1_0_INV
    );
  RXD_0_EXP_PT_1_2_INV_1053 : X_INV 
    port map (
      I => RXD_0_FBK,
      O => RXD_0_EXP_PT_1_2_INV
    );
  RXD_0_D2_PT_0_1_INV_1054 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_0_D2_PT_0_1_INV
    );
  RXD_0_D2_PT_0_3_INV_1055 : X_INV 
    port map (
      I => RXD_0_FBK,
      O => RXD_0_D2_PT_0_3_INV
    );
  RXD_0_D2_PT_1_1_INV_1056 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_0_D2_PT_1_1_INV
    );
  RXD_0_D2_PT_1_2_INV_1057 : X_INV 
    port map (
      I => UAR1_BYTE_OUT(0),
      O => RXD_0_D2_PT_1_2_INV
    );
  UAR1_BYTE_OUT_0_D2_PT_0_0_INV_1058 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_9_FBK,
      O => UAR1_BYTE_OUT_0_D2_PT_0_0_INV
    );
  CM_PANIC_ON_D2_PT_4_0_INV_1059 : X_INV 
    port map (
      I => RXD_READY_FBK,
      O => CM_PANIC_ON_D2_PT_4_0_INV
    );
  CM_PANIC_ON_D2_PT_4_1_INV_1060 : X_INV 
    port map (
      I => RXD_READY_FBK,
      O => CM_PANIC_ON_D2_PT_4_1_INV
    );
  CM_PANIC_ON_D2_PT_5_1_INV_1061 : X_INV 
    port map (
      I => RXD_4_FBK,
      O => CM_PANIC_ON_D2_PT_5_1_INV
    );
  CM_PANIC_ON_D2_PT_6_0_INV_1062 : X_INV 
    port map (
      I => RC_ADDRESS_C(0),
      O => CM_PANIC_ON_D2_PT_6_0_INV
    );
  CM_PANIC_ON_XOR_0_INV_1063 : X_INV 
    port map (
      I => CM_PANIC_ON_D1,
      O => CM_PANIC_ON_XOR_0_INV
    );
  EXP17_EXP_PT_0_1_INV_1064 : X_INV 
    port map (
      I => RXD_5_FBK,
      O => EXP17_EXP_PT_0_1_INV
    );
  EXP17_EXP_PT_1_0_INV_1065 : X_INV 
    port map (
      I => RC_ADDRESS_C(1),
      O => EXP17_EXP_PT_1_0_INV
    );
  EXP17_EXP_PT_2_1_INV_1066 : X_INV 
    port map (
      I => RXD_6_FBK,
      O => EXP17_EXP_PT_2_1_INV
    );
  EXP17_EXP_PT_3_0_INV_1067 : X_INV 
    port map (
      I => RC_ADDRESS_C(2),
      O => EXP17_EXP_PT_3_0_INV
    );
  EXP17_EXP_PT_4_1_INV_1068 : X_INV 
    port map (
      I => RXD_7_FBK,
      O => EXP17_EXP_PT_4_1_INV
    );
  EXP18_EXP_PT_2_0_INV_1069 : X_INV 
    port map (
      I => RXD_3_FBK,
      O => EXP18_EXP_PT_2_0_INV
    );
  EXP18_EXP_PT_2_1_INV_1070 : X_INV 
    port map (
      I => CM_PANIC_ON_FBK,
      O => EXP18_EXP_PT_2_1_INV
    );
  EXP18_EXP_PT_3_1_INV_1071 : X_INV 
    port map (
      I => CM_PANIC_ON_FBK,
      O => EXP18_EXP_PT_3_1_INV
    );
  EXP18_EXP_PT_4_0_INV_1072 : X_INV 
    port map (
      I => CM_PANIC_ON_FBK,
      O => EXP18_EXP_PT_4_0_INV
    );
  EXP18_EXP_PT_5_0_INV_1073 : X_INV 
    port map (
      I => RC_ADDRESS_C(3),
      O => EXP18_EXP_PT_5_0_INV
    );
  RXD_4_D2_PT_0_1_INV_1074 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_4_D2_PT_0_1_INV
    );
  RXD_4_D2_PT_0_3_INV_1075 : X_INV 
    port map (
      I => UAR1_BYTE_OUT(4),
      O => RXD_4_D2_PT_0_3_INV
    );
  RXD_4_D2_PT_1_1_INV_1076 : X_INV 
    port map (
      I => RXD_ACK,
      O => RXD_4_D2_PT_1_1_INV
    );
  RXD_4_D2_PT_1_2_INV_1077 : X_INV 
    port map (
      I => RXD_4_FBK,
      O => RXD_4_D2_PT_1_2_INV
    );
  UAR1_BYTE_OUT_4_D2_PT_0_0_INV_1078 : X_INV 
    port map (
      I => UAR1_BC1_CURRENT_STATE_5_FBK,
      O => UAR1_BYTE_OUT_4_D2_PT_0_0_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_1_0_INV_1079 : X_INV 
    port map (
      I => CM_FADE_DOWN,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_1_0_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_1_1_INV_1080 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D2_PT_1_1_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_XOR_0_INV_1081 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_D1,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_XOR_0_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_0_INV_1082 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_0_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_2_INV_1083 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_2_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_3_INV_1084 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_3_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_4_INV_1085 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_4_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_5_INV_1086 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_5_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_6_INV_1087 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_6_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_7_INV_1088 : X_INV 
    port map (
      I => FC1_CNT_6_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_7_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_8_INV_1089 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_0_8_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_0_INV_1090 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_0_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_1_INV_1091 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_1_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_2_INV_1092 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_2_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_3_INV_1093 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_3_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_4_INV_1094 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_4_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_5_INV_1095 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_5_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_6_INV_1096 : X_INV 
    port map (
      I => FC1_CNT_6_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_6_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_7_INV_1097 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_1_7_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_1_INV_1098 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_1_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_9_INV_1099 : X_INV 
    port map (
      I => LIGHT_VALUE(3),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_9_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_10_INV_1100 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_2_10_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_1_INV_1101 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_1_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_9_INV_1102 : X_INV 
    port map (
      I => LIGHT_VALUE(1),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_9_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_10_INV_1103 : X_INV 
    port map (
      I => LIGHT_VALUE(2),
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_10_INV
    );
  DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_11_INV_1104 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_EXP_PT_3_11_INV
    );
  FC1_CNT_3_RSTF_PT_0_0_INV_1105 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_3_RSTF_PT_0_0_INV
    );
  FC1_CNT_3_RSTF_PT_0_1_INV_1106 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_3_RSTF_PT_0_1_INV
    );
  FC1_CNT_3_D2_PT_2_0_INV_1107 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_3_D2_PT_2_0_INV
    );
  FC1_CNT_3_D2_PT_2_1_INV_1108 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => FC1_CNT_3_D2_PT_2_1_INV
    );
  FC1_CNT_3_D2_PT_2_2_INV_1109 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => FC1_CNT_3_D2_PT_2_2_INV
    );
  FC1_CNT_3_D2_PT_2_3_INV_1110 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => FC1_CNT_3_D2_PT_2_3_INV
    );
  FC1_CNT_3_D2_PT_2_4_INV_1111 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => FC1_CNT_3_D2_PT_2_4_INV
    );
  FC1_CNT_3_D2_PT_2_5_INV_1112 : X_INV 
    port map (
      I => FC1_CNT_6_FBK,
      O => FC1_CNT_3_D2_PT_2_5_INV
    );
  FC1_CNT_3_D2_PT_2_6_INV_1113 : X_INV 
    port map (
      I => LIGHT_VALUE(5),
      O => FC1_CNT_3_D2_PT_2_6_INV
    );
  FC1_CNT_3_D2_PT_2_7_INV_1114 : X_INV 
    port map (
      I => LIGHT_VALUE(3),
      O => FC1_CNT_3_D2_PT_2_7_INV
    );
  FC1_CNT_3_D2_PT_2_8_INV_1115 : X_INV 
    port map (
      I => LIGHT_VALUE(1),
      O => FC1_CNT_3_D2_PT_2_8_INV
    );
  FC1_CNT_3_D2_PT_2_9_INV_1116 : X_INV 
    port map (
      I => LIGHT_VALUE(2),
      O => FC1_CNT_3_D2_PT_2_9_INV
    );
  FC1_CNT_3_D2_PT_2_10_INV_1117 : X_INV 
    port map (
      I => LIGHT_VALUE(0),
      O => FC1_CNT_3_D2_PT_2_10_INV
    );
  FC1_CNT_3_D2_PT_2_11_INV_1118 : X_INV 
    port map (
      I => FC1_CNT_7_FBK,
      O => FC1_CNT_3_D2_PT_2_11_INV
    );
  FC1_CNT_3_XOR_0_INV_1119 : X_INV 
    port map (
      I => FC1_CNT_3_D1,
      O => FC1_CNT_3_XOR_0_INV
    );
  FC1_CNT_3_EXP_PT_0_0_INV_1120 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_3_EXP_PT_0_0_INV
    );
  FC1_CNT_3_EXP_PT_0_1_INV_1121 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => FC1_CNT_3_EXP_PT_0_1_INV
    );
  FC1_CNT_3_EXP_PT_0_2_INV_1122 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => FC1_CNT_3_EXP_PT_0_2_INV
    );
  FC1_CNT_3_EXP_PT_0_3_INV_1123 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => FC1_CNT_3_EXP_PT_0_3_INV
    );
  FC1_CNT_3_EXP_PT_0_4_INV_1124 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => FC1_CNT_3_EXP_PT_0_4_INV
    );
  FC1_CNT_3_EXP_PT_0_5_INV_1125 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => FC1_CNT_3_EXP_PT_0_5_INV
    );
  FC1_CNT_3_EXP_PT_0_6_INV_1126 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => FC1_CNT_3_EXP_PT_0_6_INV
    );
  FC1_CNT_3_EXP_PT_1_0_INV_1127 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_3_EXP_PT_1_0_INV
    );
  FC1_CNT_3_EXP_PT_1_1_INV_1128 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => FC1_CNT_3_EXP_PT_1_1_INV
    );
  FC1_CNT_3_EXP_PT_1_2_INV_1129 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => FC1_CNT_3_EXP_PT_1_2_INV
    );
  FC1_CNT_3_EXP_PT_1_3_INV_1130 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => FC1_CNT_3_EXP_PT_1_3_INV
    );
  FC1_CNT_3_EXP_PT_1_4_INV_1131 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => FC1_CNT_3_EXP_PT_1_4_INV
    );
  FC1_CNT_3_EXP_PT_1_5_INV_1132 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => FC1_CNT_3_EXP_PT_1_5_INV
    );
  FC1_CNT_3_EXP_PT_1_6_INV_1133 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => FC1_CNT_3_EXP_PT_1_6_INV
    );
  EXP4_EXP_PT_2_0_INV_1134 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP4_EXP_PT_2_0_INV
    );
  EXP4_EXP_PT_3_1_INV_1135 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP4_EXP_PT_3_1_INV
    );
  FC1_CNT_7_RSTF_PT_0_0_INV_1136 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_7_RSTF_PT_0_0_INV
    );
  FC1_CNT_7_RSTF_PT_0_1_INV_1137 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_7_RSTF_PT_0_1_INV
    );
  FC1_CNT_7_D2_PT_1_8_INV_1138 : X_INV 
    port map (
      I => LIGHT_VALUE(5),
      O => FC1_CNT_7_D2_PT_1_8_INV
    );
  FC1_CNT_7_D2_PT_1_9_INV_1139 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_7_D2_PT_1_9_INV
    );
  FC1_CNT_7_EXP_PT_0_1_INV_1140 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => FC1_CNT_7_EXP_PT_0_1_INV
    );
  FC1_CNT_7_EXP_PT_1_0_INV_1141 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_7_EXP_PT_1_0_INV
    );
  FC1_CNT_7_EXP_PT_1_1_INV_1142 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_7_EXP_PT_1_1_INV
    );
  FC1_CNT_7_EXP_PT_2_0_INV_1143 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => FC1_CNT_7_EXP_PT_2_0_INV
    );
  EXP3_EXP_PT_1_0_INV_1144 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP3_EXP_PT_1_0_INV
    );
  EXP3_EXP_PT_1_1_INV_1145 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP3_EXP_PT_1_1_INV
    );
  EXP3_EXP_PT_1_2_INV_1146 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP3_EXP_PT_1_2_INV
    );
  EXP3_EXP_PT_1_3_INV_1147 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP3_EXP_PT_1_3_INV
    );
  EXP3_EXP_PT_1_4_INV_1148 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP3_EXP_PT_1_4_INV
    );
  EXP3_EXP_PT_1_5_INV_1149 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => EXP3_EXP_PT_1_5_INV
    );
  EXP3_EXP_PT_1_6_INV_1150 : X_INV 
    port map (
      I => FC1_CNT_6_FBK,
      O => EXP3_EXP_PT_1_6_INV
    );
  EXP3_EXP_PT_1_7_INV_1151 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP3_EXP_PT_1_7_INV
    );
  EXP3_EXP_PT_2_0_INV_1152 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP3_EXP_PT_2_0_INV
    );
  EXP3_EXP_PT_2_1_INV_1153 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP3_EXP_PT_2_1_INV
    );
  EXP3_EXP_PT_2_2_INV_1154 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP3_EXP_PT_2_2_INV
    );
  EXP3_EXP_PT_2_3_INV_1155 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP3_EXP_PT_2_3_INV
    );
  EXP3_EXP_PT_2_4_INV_1156 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP3_EXP_PT_2_4_INV
    );
  EXP3_EXP_PT_2_5_INV_1157 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => EXP3_EXP_PT_2_5_INV
    );
  EXP3_EXP_PT_2_6_INV_1158 : X_INV 
    port map (
      I => FC1_CNT_6_FBK,
      O => EXP3_EXP_PT_2_6_INV
    );
  EXP3_EXP_PT_2_7_INV_1159 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP3_EXP_PT_2_7_INV
    );
  EXP3_EXP_PT_3_0_INV_1160 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP3_EXP_PT_3_0_INV
    );
  EXP3_EXP_PT_3_1_INV_1161 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP3_EXP_PT_3_1_INV
    );
  EXP3_EXP_PT_3_2_INV_1162 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP3_EXP_PT_3_2_INV
    );
  EXP3_EXP_PT_3_3_INV_1163 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP3_EXP_PT_3_3_INV
    );
  EXP3_EXP_PT_3_4_INV_1164 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP3_EXP_PT_3_4_INV
    );
  EXP3_EXP_PT_3_5_INV_1165 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => EXP3_EXP_PT_3_5_INV
    );
  EXP3_EXP_PT_3_6_INV_1166 : X_INV 
    port map (
      I => FC1_CNT_6_FBK,
      O => EXP3_EXP_PT_3_6_INV
    );
  EXP3_EXP_PT_3_7_INV_1167 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP3_EXP_PT_3_7_INV
    );
  EXP3_EXP_PT_4_0_INV_1168 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP3_EXP_PT_4_0_INV
    );
  EXP3_EXP_PT_4_1_INV_1169 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP3_EXP_PT_4_1_INV
    );
  EXP3_EXP_PT_4_2_INV_1170 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP3_EXP_PT_4_2_INV
    );
  EXP3_EXP_PT_4_3_INV_1171 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP3_EXP_PT_4_3_INV
    );
  EXP3_EXP_PT_4_4_INV_1172 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP3_EXP_PT_4_4_INV
    );
  EXP3_EXP_PT_4_5_INV_1173 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => EXP3_EXP_PT_4_5_INV
    );
  EXP3_EXP_PT_4_6_INV_1174 : X_INV 
    port map (
      I => FC1_CNT_6_FBK,
      O => EXP3_EXP_PT_4_6_INV
    );
  EXP3_EXP_PT_4_7_INV_1175 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP3_EXP_PT_4_7_INV
    );
  EXP3_EXP_PT_5_0_INV_1176 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP3_EXP_PT_5_0_INV
    );
  EXP3_EXP_PT_5_1_INV_1177 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP3_EXP_PT_5_1_INV
    );
  EXP3_EXP_PT_5_2_INV_1178 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP3_EXP_PT_5_2_INV
    );
  EXP3_EXP_PT_5_3_INV_1179 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP3_EXP_PT_5_3_INV
    );
  EXP3_EXP_PT_5_4_INV_1180 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP3_EXP_PT_5_4_INV
    );
  EXP3_EXP_PT_5_5_INV_1181 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => EXP3_EXP_PT_5_5_INV
    );
  EXP3_EXP_PT_5_6_INV_1182 : X_INV 
    port map (
      I => FC1_CNT_6_FBK,
      O => EXP3_EXP_PT_5_6_INV
    );
  EXP3_EXP_PT_5_7_INV_1183 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP3_EXP_PT_5_7_INV
    );
  FC1_CNT_1_RSTF_PT_0_0_INV_1184 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => FC1_CNT_1_RSTF_PT_0_0_INV
    );
  FC1_CNT_1_RSTF_PT_0_1_INV_1185 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => FC1_CNT_1_RSTF_PT_0_1_INV
    );
  FC1_CNT_1_D2_PT_4_0_INV_1186 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => FC1_CNT_1_D2_PT_4_0_INV
    );
  FC1_CNT_1_D2_PT_4_1_INV_1187 : X_INV 
    port map (
      I => LIGHT_VALUE_5_FBK,
      O => FC1_CNT_1_D2_PT_4_1_INV
    );
  FC1_CNT_1_D2_PT_4_2_INV_1188 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => FC1_CNT_1_D2_PT_4_2_INV
    );
  FC1_CNT_1_D2_PT_4_3_INV_1189 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => FC1_CNT_1_D2_PT_4_3_INV
    );
  FC1_CNT_1_D2_PT_4_4_INV_1190 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => FC1_CNT_1_D2_PT_4_4_INV
    );
  FC1_CNT_1_D2_PT_4_5_INV_1191 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => FC1_CNT_1_D2_PT_4_5_INV
    );
  FC1_CNT_1_D2_PT_4_6_INV_1192 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => FC1_CNT_1_D2_PT_4_6_INV
    );
  FC1_CNT_1_D2_PT_4_7_INV_1193 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => FC1_CNT_1_D2_PT_4_7_INV
    );
  FC1_CNT_1_D2_PT_4_8_INV_1194 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => FC1_CNT_1_D2_PT_4_8_INV
    );
  FC1_CNT_1_D2_PT_4_9_INV_1195 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => FC1_CNT_1_D2_PT_4_9_INV
    );
  FC1_CNT_1_D2_PT_4_10_INV_1196 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => FC1_CNT_1_D2_PT_4_10_INV
    );
  FC1_CNT_1_D2_PT_4_11_INV_1197 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => FC1_CNT_1_D2_PT_4_11_INV
    );
  FC1_CNT_1_D2_PT_4_12_INV_1198 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => FC1_CNT_1_D2_PT_4_12_INV
    );
  FC1_CNT_1_D2_PT_4_13_INV_1199 : X_INV 
    port map (
      I => LIGHT_VALUE(4),
      O => FC1_CNT_1_D2_PT_4_13_INV
    );
  FC1_CNT_1_XOR_0_INV_1200 : X_INV 
    port map (
      I => FC1_CNT_1_D1,
      O => FC1_CNT_1_XOR_0_INV
    );
  FC1_CNT_0_RSTF_PT_0_0_INV_1201 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => FC1_CNT_0_RSTF_PT_0_0_INV
    );
  FC1_CNT_0_RSTF_PT_0_1_INV_1202 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => FC1_CNT_0_RSTF_PT_0_1_INV
    );
  FC1_CNT_0_XOR_0_INV_1203 : X_INV 
    port map (
      I => FC1_CNT_0_D1,
      O => FC1_CNT_0_XOR_0_INV
    );
  FC1_CNT_0_EXP_PT_1_0_INV_1204 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => FC1_CNT_0_EXP_PT_1_0_INV
    );
  FC1_CNT_0_EXP_PT_1_1_INV_1205 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => FC1_CNT_0_EXP_PT_1_1_INV
    );
  FC1_CNT_0_EXP_PT_2_0_INV_1206 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => FC1_CNT_0_EXP_PT_2_0_INV
    );
  EXP12_EXP_PT_0_0_INV_1207 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => EXP12_EXP_PT_0_0_INV
    );
  EXP12_EXP_PT_0_1_INV_1208 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => EXP12_EXP_PT_0_1_INV
    );
  EXP12_EXP_PT_1_0_INV_1209 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => EXP12_EXP_PT_1_0_INV
    );
  EXP12_EXP_PT_2_0_INV_1210 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => EXP12_EXP_PT_2_0_INV
    );
  EXP12_EXP_PT_3_0_INV_1211 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => EXP12_EXP_PT_3_0_INV
    );
  EXP12_EXP_PT_4_1_INV_1212 : X_INV 
    port map (
      I => LIGHT_VALUE_5_FBK,
      O => EXP12_EXP_PT_4_1_INV
    );
  EXP12_EXP_PT_4_2_INV_1213 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => EXP12_EXP_PT_4_2_INV
    );
  EXP12_EXP_PT_4_3_INV_1214 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => EXP12_EXP_PT_4_3_INV
    );
  EXP12_EXP_PT_4_4_INV_1215 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => EXP12_EXP_PT_4_4_INV
    );
  EXP12_EXP_PT_4_5_INV_1216 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => EXP12_EXP_PT_4_5_INV
    );
  EXP12_EXP_PT_4_6_INV_1217 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => EXP12_EXP_PT_4_6_INV
    );
  EXP12_EXP_PT_4_7_INV_1218 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => EXP12_EXP_PT_4_7_INV
    );
  EXP12_EXP_PT_4_8_INV_1219 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => EXP12_EXP_PT_4_8_INV
    );
  EXP12_EXP_PT_4_9_INV_1220 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => EXP12_EXP_PT_4_9_INV
    );
  EXP12_EXP_PT_4_10_INV_1221 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => EXP12_EXP_PT_4_10_INV
    );
  EXP12_EXP_PT_4_11_INV_1222 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => EXP12_EXP_PT_4_11_INV
    );
  EXP12_EXP_PT_4_12_INV_1223 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => EXP12_EXP_PT_4_12_INV
    );
  EXP12_EXP_PT_4_13_INV_1224 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => EXP12_EXP_PT_4_13_INV
    );
  EXP12_EXP_PT_4_14_INV_1225 : X_INV 
    port map (
      I => LIGHT_VALUE(4),
      O => EXP12_EXP_PT_4_14_INV
    );
  LIGHT_VALUE_5_SETF_PT_0_0_INV_1226 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => LIGHT_VALUE_5_SETF_PT_0_0_INV
    );
  LIGHT_VALUE_5_SETF_PT_0_1_INV_1227 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_5_SETF_PT_0_1_INV
    );
  LIGHT_VALUE_5_D2_PT_1_0_INV_1228 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => LIGHT_VALUE_5_D2_PT_1_0_INV
    );
  LIGHT_VALUE_5_D2_PT_1_2_INV_1229 : X_INV 
    port map (
      I => LIGHT_VALUE_5_FBK,
      O => LIGHT_VALUE_5_D2_PT_1_2_INV
    );
  LIGHT_VALUE_5_EXP_PT_0_1_INV_1230 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_5_EXP_PT_0_1_INV
    );
  LIGHT_VALUE_5_EXP_PT_0_3_INV_1231 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_5_EXP_PT_0_3_INV
    );
  LIGHT_VALUE_5_EXP_PT_0_4_INV_1232 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => LIGHT_VALUE_5_EXP_PT_0_4_INV
    );
  LIGHT_VALUE_5_EXP_PT_0_5_INV_1233 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => LIGHT_VALUE_5_EXP_PT_0_5_INV
    );
  LIGHT_VALUE_5_EXP_PT_0_6_INV_1234 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => LIGHT_VALUE_5_EXP_PT_0_6_INV
    );
  LIGHT_VALUE_5_EXP_PT_0_7_INV_1235 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => LIGHT_VALUE_5_EXP_PT_0_7_INV
    );
  LIGHT_VALUE_5_EXP_PT_0_8_INV_1236 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => LIGHT_VALUE_5_EXP_PT_0_8_INV
    );
  LIGHT_VALUE_5_EXP_PT_0_9_INV_1237 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => LIGHT_VALUE_5_EXP_PT_0_9_INV
    );
  LIGHT_VALUE_5_EXP_PT_0_10_INV_1238 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => LIGHT_VALUE_5_EXP_PT_0_10_INV
    );
  LIGHT_VALUE_5_EXP_PT_0_11_INV_1239 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => LIGHT_VALUE_5_EXP_PT_0_11_INV
    );
  LIGHT_VALUE_5_EXP_PT_0_12_INV_1240 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => LIGHT_VALUE_5_EXP_PT_0_12_INV
    );
  LIGHT_VALUE_5_EXP_PT_0_13_INV_1241 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => LIGHT_VALUE_5_EXP_PT_0_13_INV
    );
  LIGHT_VALUE_5_EXP_PT_1_1_INV_1242 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_5_EXP_PT_1_1_INV
    );
  LIGHT_VALUE_5_EXP_PT_1_2_INV_1243 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_5_EXP_PT_1_2_INV
    );
  LIGHT_VALUE_5_EXP_PT_1_3_INV_1244 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => LIGHT_VALUE_5_EXP_PT_1_3_INV
    );
  LIGHT_VALUE_5_EXP_PT_1_4_INV_1245 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => LIGHT_VALUE_5_EXP_PT_1_4_INV
    );
  LIGHT_VALUE_5_EXP_PT_1_5_INV_1246 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => LIGHT_VALUE_5_EXP_PT_1_5_INV
    );
  LIGHT_VALUE_5_EXP_PT_1_6_INV_1247 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => LIGHT_VALUE_5_EXP_PT_1_6_INV
    );
  LIGHT_VALUE_5_EXP_PT_1_7_INV_1248 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => LIGHT_VALUE_5_EXP_PT_1_7_INV
    );
  LIGHT_VALUE_5_EXP_PT_1_8_INV_1249 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => LIGHT_VALUE_5_EXP_PT_1_8_INV
    );
  LIGHT_VALUE_5_EXP_PT_1_9_INV_1250 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => LIGHT_VALUE_5_EXP_PT_1_9_INV
    );
  LIGHT_VALUE_5_EXP_PT_1_10_INV_1251 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => LIGHT_VALUE_5_EXP_PT_1_10_INV
    );
  LIGHT_VALUE_5_EXP_PT_1_11_INV_1252 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => LIGHT_VALUE_5_EXP_PT_1_11_INV
    );
  LIGHT_VALUE_5_EXP_PT_1_12_INV_1253 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => LIGHT_VALUE_5_EXP_PT_1_12_INV
    );
  LIGHT_VALUE_5_EXP_PT_2_0_INV_1254 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => LIGHT_VALUE_5_EXP_PT_2_0_INV
    );
  LIGHT_VALUE_5_EXP_PT_2_13_INV_1255 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => LIGHT_VALUE_5_EXP_PT_2_13_INV
    );
  LIGHT_VALUE_5_EXP_PT_2_14_INV_1256 : X_INV 
    port map (
      I => LIGHT_VALUE(4),
      O => LIGHT_VALUE_5_EXP_PT_2_14_INV
    );
  TD1_CNT_0_RSTF_PT_0_0_INV_1257 : X_INV 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM,
      O => TD1_CNT_0_RSTF_PT_0_0_INV
    );
  TD1_CNT_0_RSTF_PT_0_1_INV_1258 : X_INV 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM,
      O => TD1_CNT_0_RSTF_PT_0_1_INV
    );
  TD1_CNT_0_D2_PT_0_0_INV_1259 : X_INV 
    port map (
      I => TD1_CNT_0_FBK,
      O => TD1_CNT_0_D2_PT_0_0_INV
    );
  TD1_CNT_0_D2_PT_0_1_INV_1260 : X_INV 
    port map (
      I => TD1_CNT_0_FBK,
      O => TD1_CNT_0_D2_PT_0_1_INV
    );
  TD1_CNT_0_EXP_PT_0_1_INV_1261 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => TD1_CNT_0_EXP_PT_0_1_INV
    );
  TD1_CNT_0_EXP_PT_0_3_INV_1262 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => TD1_CNT_0_EXP_PT_0_3_INV
    );
  TD1_CNT_0_EXP_PT_0_4_INV_1263 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => TD1_CNT_0_EXP_PT_0_4_INV
    );
  TD1_CNT_0_EXP_PT_0_5_INV_1264 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => TD1_CNT_0_EXP_PT_0_5_INV
    );
  TD1_CNT_0_EXP_PT_0_6_INV_1265 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => TD1_CNT_0_EXP_PT_0_6_INV
    );
  TD1_CNT_0_EXP_PT_0_7_INV_1266 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => TD1_CNT_0_EXP_PT_0_7_INV
    );
  TD1_CNT_0_EXP_PT_0_8_INV_1267 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => TD1_CNT_0_EXP_PT_0_8_INV
    );
  TD1_CNT_0_EXP_PT_0_9_INV_1268 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => TD1_CNT_0_EXP_PT_0_9_INV
    );
  TD1_CNT_0_EXP_PT_0_10_INV_1269 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => TD1_CNT_0_EXP_PT_0_10_INV
    );
  TD1_CNT_0_EXP_PT_0_11_INV_1270 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => TD1_CNT_0_EXP_PT_0_11_INV
    );
  TD1_CNT_0_EXP_PT_0_12_INV_1271 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => TD1_CNT_0_EXP_PT_0_12_INV
    );
  TD1_CNT_0_EXP_PT_0_13_INV_1272 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => TD1_CNT_0_EXP_PT_0_13_INV
    );
  TD1_CNT_0_EXP_PT_0_14_INV_1273 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => TD1_CNT_0_EXP_PT_0_14_INV
    );
  TD1_CNT_0_EXP_PT_0_15_INV_1274 : X_INV 
    port map (
      I => LIGHT_VALUE(4),
      O => TD1_CNT_0_EXP_PT_0_15_INV
    );
  TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0_0_INV_1275 : X_INV 
    port map (
      I => RESET_C,
      O => TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0_0_INV
    );
  TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0_1_INV_1276 : X_INV 
    port map (
      I => ZERO_DETECT_C,
      O => TD1_CNT_5_TD1_CNT_5_SETF_INT_D2_PT_0_1_INV
    );
  FC1_CNT_2_RSTF_PT_0_0_INV_1277 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => FC1_CNT_2_RSTF_PT_0_0_INV
    );
  FC1_CNT_2_RSTF_PT_0_1_INV_1278 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => FC1_CNT_2_RSTF_PT_0_1_INV
    );
  FC1_CNT_2_D2_PT_2_0_INV_1279 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => FC1_CNT_2_D2_PT_2_0_INV
    );
  FC1_CNT_2_D2_PT_2_1_INV_1280 : X_INV 
    port map (
      I => LIGHT_VALUE_5_FBK,
      O => FC1_CNT_2_D2_PT_2_1_INV
    );
  FC1_CNT_2_D2_PT_2_2_INV_1281 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => FC1_CNT_2_D2_PT_2_2_INV
    );
  FC1_CNT_2_D2_PT_2_3_INV_1282 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => FC1_CNT_2_D2_PT_2_3_INV
    );
  FC1_CNT_2_D2_PT_2_4_INV_1283 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => FC1_CNT_2_D2_PT_2_4_INV
    );
  FC1_CNT_2_D2_PT_2_5_INV_1284 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => FC1_CNT_2_D2_PT_2_5_INV
    );
  FC1_CNT_2_D2_PT_2_6_INV_1285 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => FC1_CNT_2_D2_PT_2_6_INV
    );
  FC1_CNT_2_D2_PT_2_7_INV_1286 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => FC1_CNT_2_D2_PT_2_7_INV
    );
  FC1_CNT_2_D2_PT_2_8_INV_1287 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => FC1_CNT_2_D2_PT_2_8_INV
    );
  FC1_CNT_2_D2_PT_2_9_INV_1288 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => FC1_CNT_2_D2_PT_2_9_INV
    );
  FC1_CNT_2_D2_PT_2_10_INV_1289 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => FC1_CNT_2_D2_PT_2_10_INV
    );
  FC1_CNT_2_D2_PT_2_11_INV_1290 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => FC1_CNT_2_D2_PT_2_11_INV
    );
  FC1_CNT_2_D2_PT_2_12_INV_1291 : X_INV 
    port map (
      I => LIGHT_VALUE(4),
      O => FC1_CNT_2_D2_PT_2_12_INV
    );
  FC1_CNT_2_XOR_0_INV_1292 : X_INV 
    port map (
      I => FC1_CNT_2_D1,
      O => FC1_CNT_2_XOR_0_INV
    );
  FC1_CNT_2_EXP_PT_0_1_INV_1293 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => FC1_CNT_2_EXP_PT_0_1_INV
    );
  FC1_CNT_2_EXP_PT_0_2_INV_1294 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => FC1_CNT_2_EXP_PT_0_2_INV
    );
  FC1_CNT_2_EXP_PT_0_3_INV_1295 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => FC1_CNT_2_EXP_PT_0_3_INV
    );
  FC1_CNT_2_EXP_PT_0_4_INV_1296 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => FC1_CNT_2_EXP_PT_0_4_INV
    );
  FC1_CNT_2_EXP_PT_0_5_INV_1297 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => FC1_CNT_2_EXP_PT_0_5_INV
    );
  FC1_CNT_2_EXP_PT_0_6_INV_1298 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => FC1_CNT_2_EXP_PT_0_6_INV
    );
  FC1_CNT_2_EXP_PT_0_7_INV_1299 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => FC1_CNT_2_EXP_PT_0_7_INV
    );
  FC1_CNT_2_EXP_PT_0_8_INV_1300 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => FC1_CNT_2_EXP_PT_0_8_INV
    );
  FC1_CNT_2_EXP_PT_0_9_INV_1301 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => FC1_CNT_2_EXP_PT_0_9_INV
    );
  FC1_CNT_2_EXP_PT_1_1_INV_1302 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => FC1_CNT_2_EXP_PT_1_1_INV
    );
  FC1_CNT_2_EXP_PT_1_2_INV_1303 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => FC1_CNT_2_EXP_PT_1_2_INV
    );
  FC1_CNT_2_EXP_PT_1_3_INV_1304 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => FC1_CNT_2_EXP_PT_1_3_INV
    );
  FC1_CNT_2_EXP_PT_1_4_INV_1305 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => FC1_CNT_2_EXP_PT_1_4_INV
    );
  FC1_CNT_2_EXP_PT_1_5_INV_1306 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => FC1_CNT_2_EXP_PT_1_5_INV
    );
  FC1_CNT_2_EXP_PT_1_6_INV_1307 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => FC1_CNT_2_EXP_PT_1_6_INV
    );
  FC1_CNT_2_EXP_PT_1_7_INV_1308 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => FC1_CNT_2_EXP_PT_1_7_INV
    );
  FC1_CNT_2_EXP_PT_1_8_INV_1309 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => FC1_CNT_2_EXP_PT_1_8_INV
    );
  FC1_CNT_2_EXP_PT_1_9_INV_1310 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => FC1_CNT_2_EXP_PT_1_9_INV
    );
  EXP14_EXP_PT_2_0_INV_1311 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => EXP14_EXP_PT_2_0_INV
    );
  EXP14_EXP_PT_2_1_INV_1312 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => EXP14_EXP_PT_2_1_INV
    );
  EXP14_EXP_PT_3_1_INV_1313 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => EXP14_EXP_PT_3_1_INV
    );
  LIGHT_VALUE_1_SETF_PT_0_0_INV_1314 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => LIGHT_VALUE_1_SETF_PT_0_0_INV
    );
  LIGHT_VALUE_1_SETF_PT_0_1_INV_1315 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_1_SETF_PT_0_1_INV
    );
  LIGHT_VALUE_1_D2_PT_1_1_INV_1316 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_1_D2_PT_1_1_INV
    );
  LIGHT_VALUE_1_D2_PT_1_2_INV_1317 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_1_D2_PT_1_2_INV
    );
  LIGHT_VALUE_1_D2_PT_1_3_INV_1318 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => LIGHT_VALUE_1_D2_PT_1_3_INV
    );
  LIGHT_VALUE_1_D2_PT_1_4_INV_1319 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => LIGHT_VALUE_1_D2_PT_1_4_INV
    );
  LIGHT_VALUE_1_D2_PT_1_5_INV_1320 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => LIGHT_VALUE_1_D2_PT_1_5_INV
    );
  LIGHT_VALUE_1_D2_PT_1_6_INV_1321 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => LIGHT_VALUE_1_D2_PT_1_6_INV
    );
  LIGHT_VALUE_1_D2_PT_1_7_INV_1322 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => LIGHT_VALUE_1_D2_PT_1_7_INV
    );
  LIGHT_VALUE_1_D2_PT_1_8_INV_1323 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => LIGHT_VALUE_1_D2_PT_1_8_INV
    );
  LIGHT_VALUE_1_D2_PT_1_9_INV_1324 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => LIGHT_VALUE_1_D2_PT_1_9_INV
    );
  LIGHT_VALUE_1_D2_PT_1_11_INV_1325 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => LIGHT_VALUE_1_D2_PT_1_11_INV
    );
  LIGHT_VALUE_1_D2_PT_2_1_INV_1326 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_1_D2_PT_2_1_INV
    );
  LIGHT_VALUE_1_D2_PT_2_2_INV_1327 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_1_D2_PT_2_2_INV
    );
  LIGHT_VALUE_1_D2_PT_2_3_INV_1328 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => LIGHT_VALUE_1_D2_PT_2_3_INV
    );
  LIGHT_VALUE_1_D2_PT_2_4_INV_1329 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => LIGHT_VALUE_1_D2_PT_2_4_INV
    );
  LIGHT_VALUE_1_D2_PT_2_5_INV_1330 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => LIGHT_VALUE_1_D2_PT_2_5_INV
    );
  LIGHT_VALUE_1_D2_PT_2_6_INV_1331 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => LIGHT_VALUE_1_D2_PT_2_6_INV
    );
  LIGHT_VALUE_1_D2_PT_2_7_INV_1332 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => LIGHT_VALUE_1_D2_PT_2_7_INV
    );
  LIGHT_VALUE_1_D2_PT_2_8_INV_1333 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => LIGHT_VALUE_1_D2_PT_2_8_INV
    );
  LIGHT_VALUE_1_D2_PT_2_9_INV_1334 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => LIGHT_VALUE_1_D2_PT_2_9_INV
    );
  LIGHT_VALUE_1_D2_PT_2_11_INV_1335 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => LIGHT_VALUE_1_D2_PT_2_11_INV
    );
  LIGHT_VALUE_1_D2_PT_3_0_INV_1336 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => LIGHT_VALUE_1_D2_PT_3_0_INV
    );
  LIGHT_VALUE_1_D2_PT_3_2_INV_1337 : X_INV 
    port map (
      I => LIGHT_VALUE_5_FBK,
      O => LIGHT_VALUE_1_D2_PT_3_2_INV
    );
  LIGHT_VALUE_1_EXP_PT_0_1_INV_1338 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_1_EXP_PT_0_1_INV
    );
  EXP13_EXP_PT_0_1_INV_1339 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => EXP13_EXP_PT_0_1_INV
    );
  EXP13_EXP_PT_0_3_INV_1340 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => EXP13_EXP_PT_0_3_INV
    );
  EXP13_EXP_PT_0_4_INV_1341 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => EXP13_EXP_PT_0_4_INV
    );
  EXP13_EXP_PT_0_5_INV_1342 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => EXP13_EXP_PT_0_5_INV
    );
  EXP13_EXP_PT_0_6_INV_1343 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => EXP13_EXP_PT_0_6_INV
    );
  EXP13_EXP_PT_0_7_INV_1344 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => EXP13_EXP_PT_0_7_INV
    );
  EXP13_EXP_PT_0_8_INV_1345 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => EXP13_EXP_PT_0_8_INV
    );
  EXP13_EXP_PT_0_9_INV_1346 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => EXP13_EXP_PT_0_9_INV
    );
  EXP13_EXP_PT_0_10_INV_1347 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => EXP13_EXP_PT_0_10_INV
    );
  EXP13_EXP_PT_0_11_INV_1348 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => EXP13_EXP_PT_0_11_INV
    );
  EXP13_EXP_PT_1_1_INV_1349 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => EXP13_EXP_PT_1_1_INV
    );
  EXP13_EXP_PT_1_2_INV_1350 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => EXP13_EXP_PT_1_2_INV
    );
  EXP13_EXP_PT_1_3_INV_1351 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => EXP13_EXP_PT_1_3_INV
    );
  EXP13_EXP_PT_1_4_INV_1352 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => EXP13_EXP_PT_1_4_INV
    );
  EXP13_EXP_PT_1_5_INV_1353 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => EXP13_EXP_PT_1_5_INV
    );
  EXP13_EXP_PT_1_6_INV_1354 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => EXP13_EXP_PT_1_6_INV
    );
  EXP13_EXP_PT_1_7_INV_1355 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => EXP13_EXP_PT_1_7_INV
    );
  EXP13_EXP_PT_1_8_INV_1356 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => EXP13_EXP_PT_1_8_INV
    );
  EXP13_EXP_PT_1_9_INV_1357 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => EXP13_EXP_PT_1_9_INV
    );
  EXP13_EXP_PT_1_10_INV_1358 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => EXP13_EXP_PT_1_10_INV
    );
  EXP13_EXP_PT_2_1_INV_1359 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => EXP13_EXP_PT_2_1_INV
    );
  EXP13_EXP_PT_2_2_INV_1360 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => EXP13_EXP_PT_2_2_INV
    );
  EXP13_EXP_PT_2_3_INV_1361 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => EXP13_EXP_PT_2_3_INV
    );
  EXP13_EXP_PT_2_4_INV_1362 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => EXP13_EXP_PT_2_4_INV
    );
  EXP13_EXP_PT_2_5_INV_1363 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => EXP13_EXP_PT_2_5_INV
    );
  EXP13_EXP_PT_2_6_INV_1364 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => EXP13_EXP_PT_2_6_INV
    );
  EXP13_EXP_PT_2_7_INV_1365 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => EXP13_EXP_PT_2_7_INV
    );
  EXP13_EXP_PT_2_8_INV_1366 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => EXP13_EXP_PT_2_8_INV
    );
  EXP13_EXP_PT_2_9_INV_1367 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => EXP13_EXP_PT_2_9_INV
    );
  EXP13_EXP_PT_2_10_INV_1368 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => EXP13_EXP_PT_2_10_INV
    );
  EXP13_EXP_PT_3_0_INV_1369 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => EXP13_EXP_PT_3_0_INV
    );
  EXP13_EXP_PT_3_11_INV_1370 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => EXP13_EXP_PT_3_11_INV
    );
  EXP13_EXP_PT_3_12_INV_1371 : X_INV 
    port map (
      I => LIGHT_VALUE(4),
      O => EXP13_EXP_PT_3_12_INV
    );
  EXP13_EXP_PT_4_0_INV_1372 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => EXP13_EXP_PT_4_0_INV
    );
  EXP13_EXP_PT_4_10_INV_1373 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => EXP13_EXP_PT_4_10_INV
    );
  EXP13_EXP_PT_4_11_INV_1374 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => EXP13_EXP_PT_4_11_INV
    );
  EXP13_EXP_PT_4_13_INV_1375 : X_INV 
    port map (
      I => LIGHT_VALUE(4),
      O => EXP13_EXP_PT_4_13_INV
    );
  FC1_CNT_4_RSTF_PT_0_0_INV_1376 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_4_RSTF_PT_0_0_INV
    );
  FC1_CNT_4_RSTF_PT_0_1_INV_1377 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_4_RSTF_PT_0_1_INV
    );
  FC1_CNT_4_D2_PT_2_5_INV_1378 : X_INV 
    port map (
      I => LIGHT_VALUE(5),
      O => FC1_CNT_4_D2_PT_2_5_INV
    );
  FC1_CNT_4_D2_PT_2_6_INV_1379 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_4_D2_PT_2_6_INV
    );
  FC1_CNT_4_D2_PT_3_0_INV_1380 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_4_D2_PT_3_0_INV
    );
  FC1_CNT_4_D2_PT_3_1_INV_1381 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => FC1_CNT_4_D2_PT_3_1_INV
    );
  FC1_CNT_4_D2_PT_3_2_INV_1382 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => FC1_CNT_4_D2_PT_3_2_INV
    );
  FC1_CNT_4_D2_PT_3_3_INV_1383 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => FC1_CNT_4_D2_PT_3_3_INV
    );
  FC1_CNT_4_D2_PT_3_5_INV_1384 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => FC1_CNT_4_D2_PT_3_5_INV
    );
  FC1_CNT_4_D2_PT_4_0_INV_1385 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_4_D2_PT_4_0_INV
    );
  FC1_CNT_4_D2_PT_4_1_INV_1386 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => FC1_CNT_4_D2_PT_4_1_INV
    );
  FC1_CNT_4_D2_PT_4_2_INV_1387 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => FC1_CNT_4_D2_PT_4_2_INV
    );
  FC1_CNT_4_D2_PT_4_3_INV_1388 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => FC1_CNT_4_D2_PT_4_3_INV
    );
  FC1_CNT_4_D2_PT_4_5_INV_1389 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => FC1_CNT_4_D2_PT_4_5_INV
    );
  FC1_CNT_4_D2_PT_5_0_INV_1390 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_4_D2_PT_5_0_INV
    );
  FC1_CNT_4_D2_PT_5_1_INV_1391 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => FC1_CNT_4_D2_PT_5_1_INV
    );
  FC1_CNT_4_D2_PT_5_2_INV_1392 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => FC1_CNT_4_D2_PT_5_2_INV
    );
  FC1_CNT_4_D2_PT_5_3_INV_1393 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => FC1_CNT_4_D2_PT_5_3_INV
    );
  FC1_CNT_4_D2_PT_5_4_INV_1394 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => FC1_CNT_4_D2_PT_5_4_INV
    );
  EXP8_EXP_PT_1_0_INV_1395 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP8_EXP_PT_1_0_INV
    );
  EXP8_EXP_PT_1_1_INV_1396 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP8_EXP_PT_1_1_INV
    );
  EXP8_EXP_PT_1_2_INV_1397 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP8_EXP_PT_1_2_INV
    );
  EXP8_EXP_PT_1_3_INV_1398 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP8_EXP_PT_1_3_INV
    );
  EXP8_EXP_PT_1_5_INV_1399 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP8_EXP_PT_1_5_INV
    );
  EXP8_EXP_PT_2_0_INV_1400 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP8_EXP_PT_2_0_INV
    );
  EXP8_EXP_PT_2_1_INV_1401 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP8_EXP_PT_2_1_INV
    );
  EXP8_EXP_PT_2_2_INV_1402 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP8_EXP_PT_2_2_INV
    );
  EXP8_EXP_PT_2_3_INV_1403 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP8_EXP_PT_2_3_INV
    );
  EXP8_EXP_PT_2_4_INV_1404 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP8_EXP_PT_2_4_INV
    );
  EXP8_EXP_PT_3_0_INV_1405 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP8_EXP_PT_3_0_INV
    );
  EXP8_EXP_PT_3_1_INV_1406 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP8_EXP_PT_3_1_INV
    );
  EXP8_EXP_PT_3_2_INV_1407 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP8_EXP_PT_3_2_INV
    );
  EXP8_EXP_PT_3_3_INV_1408 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP8_EXP_PT_3_3_INV
    );
  EXP8_EXP_PT_3_4_INV_1409 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP8_EXP_PT_3_4_INV
    );
  EXP8_EXP_PT_4_0_INV_1410 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP8_EXP_PT_4_0_INV
    );
  EXP8_EXP_PT_4_1_INV_1411 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP8_EXP_PT_4_1_INV
    );
  EXP8_EXP_PT_4_2_INV_1412 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP8_EXP_PT_4_2_INV
    );
  EXP8_EXP_PT_4_3_INV_1413 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP8_EXP_PT_4_3_INV
    );
  EXP8_EXP_PT_4_4_INV_1414 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP8_EXP_PT_4_4_INV
    );
  EXP8_EXP_PT_5_0_INV_1415 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP8_EXP_PT_5_0_INV
    );
  EXP8_EXP_PT_5_1_INV_1416 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP8_EXP_PT_5_1_INV
    );
  EXP8_EXP_PT_5_2_INV_1417 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP8_EXP_PT_5_2_INV
    );
  EXP8_EXP_PT_5_3_INV_1418 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP8_EXP_PT_5_3_INV
    );
  EXP8_EXP_PT_5_4_INV_1419 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP8_EXP_PT_5_4_INV
    );
  FC1_CNT_5_RSTF_PT_0_0_INV_1420 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_5_RSTF_PT_0_0_INV
    );
  FC1_CNT_5_RSTF_PT_0_1_INV_1421 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_5_RSTF_PT_0_1_INV
    );
  FC1_CNT_5_D2_PT_1_6_INV_1422 : X_INV 
    port map (
      I => LIGHT_VALUE(5),
      O => FC1_CNT_5_D2_PT_1_6_INV
    );
  FC1_CNT_5_D2_PT_1_7_INV_1423 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_5_D2_PT_1_7_INV
    );
  FC1_CNT_5_D2_PT_2_0_INV_1424 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_5_D2_PT_2_0_INV
    );
  FC1_CNT_5_D2_PT_2_1_INV_1425 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => FC1_CNT_5_D2_PT_2_1_INV
    );
  FC1_CNT_5_D2_PT_2_2_INV_1426 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => FC1_CNT_5_D2_PT_2_2_INV
    );
  FC1_CNT_5_D2_PT_2_3_INV_1427 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => FC1_CNT_5_D2_PT_2_3_INV
    );
  FC1_CNT_5_D2_PT_2_4_INV_1428 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => FC1_CNT_5_D2_PT_2_4_INV
    );
  FC1_CNT_5_D2_PT_2_6_INV_1429 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => FC1_CNT_5_D2_PT_2_6_INV
    );
  FC1_CNT_5_D2_PT_3_0_INV_1430 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_5_D2_PT_3_0_INV
    );
  FC1_CNT_5_D2_PT_3_1_INV_1431 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => FC1_CNT_5_D2_PT_3_1_INV
    );
  FC1_CNT_5_D2_PT_3_2_INV_1432 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => FC1_CNT_5_D2_PT_3_2_INV
    );
  FC1_CNT_5_D2_PT_3_3_INV_1433 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => FC1_CNT_5_D2_PT_3_3_INV
    );
  FC1_CNT_5_D2_PT_3_4_INV_1434 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => FC1_CNT_5_D2_PT_3_4_INV
    );
  FC1_CNT_5_D2_PT_3_5_INV_1435 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => FC1_CNT_5_D2_PT_3_5_INV
    );
  FC1_CNT_5_EXP_PT_0_1_INV_1436 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => FC1_CNT_5_EXP_PT_0_1_INV
    );
  FC1_CNT_5_EXP_PT_0_6_INV_1437 : X_INV 
    port map (
      I => LIGHT_VALUE(1),
      O => FC1_CNT_5_EXP_PT_0_6_INV
    );
  FC1_CNT_5_EXP_PT_0_7_INV_1438 : X_INV 
    port map (
      I => LIGHT_VALUE(2),
      O => FC1_CNT_5_EXP_PT_0_7_INV
    );
  FC1_CNT_5_EXP_PT_0_8_INV_1439 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_5_EXP_PT_0_8_INV
    );
  EXP7_EXP_PT_1_0_INV_1440 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP7_EXP_PT_1_0_INV
    );
  EXP7_EXP_PT_1_1_INV_1441 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP7_EXP_PT_1_1_INV
    );
  EXP7_EXP_PT_1_2_INV_1442 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP7_EXP_PT_1_2_INV
    );
  EXP7_EXP_PT_1_3_INV_1443 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP7_EXP_PT_1_3_INV
    );
  EXP7_EXP_PT_1_4_INV_1444 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP7_EXP_PT_1_4_INV
    );
  EXP7_EXP_PT_1_6_INV_1445 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP7_EXP_PT_1_6_INV
    );
  EXP7_EXP_PT_2_0_INV_1446 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP7_EXP_PT_2_0_INV
    );
  EXP7_EXP_PT_2_1_INV_1447 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP7_EXP_PT_2_1_INV
    );
  EXP7_EXP_PT_2_2_INV_1448 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP7_EXP_PT_2_2_INV
    );
  EXP7_EXP_PT_2_3_INV_1449 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP7_EXP_PT_2_3_INV
    );
  EXP7_EXP_PT_2_4_INV_1450 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP7_EXP_PT_2_4_INV
    );
  EXP7_EXP_PT_2_5_INV_1451 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP7_EXP_PT_2_5_INV
    );
  EXP7_EXP_PT_3_0_INV_1452 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP7_EXP_PT_3_0_INV
    );
  EXP7_EXP_PT_3_1_INV_1453 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP7_EXP_PT_3_1_INV
    );
  EXP7_EXP_PT_3_2_INV_1454 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP7_EXP_PT_3_2_INV
    );
  EXP7_EXP_PT_3_3_INV_1455 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP7_EXP_PT_3_3_INV
    );
  EXP7_EXP_PT_3_4_INV_1456 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP7_EXP_PT_3_4_INV
    );
  EXP7_EXP_PT_3_5_INV_1457 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP7_EXP_PT_3_5_INV
    );
  EXP7_EXP_PT_4_0_INV_1458 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP7_EXP_PT_4_0_INV
    );
  EXP7_EXP_PT_4_1_INV_1459 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP7_EXP_PT_4_1_INV
    );
  EXP7_EXP_PT_4_2_INV_1460 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP7_EXP_PT_4_2_INV
    );
  EXP7_EXP_PT_4_3_INV_1461 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP7_EXP_PT_4_3_INV
    );
  EXP7_EXP_PT_4_4_INV_1462 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP7_EXP_PT_4_4_INV
    );
  EXP7_EXP_PT_4_5_INV_1463 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP7_EXP_PT_4_5_INV
    );
  EXP7_EXP_PT_5_0_INV_1464 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP7_EXP_PT_5_0_INV
    );
  EXP7_EXP_PT_5_1_INV_1465 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP7_EXP_PT_5_1_INV
    );
  EXP7_EXP_PT_5_2_INV_1466 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP7_EXP_PT_5_2_INV
    );
  EXP7_EXP_PT_5_3_INV_1467 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP7_EXP_PT_5_3_INV
    );
  EXP7_EXP_PT_5_4_INV_1468 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP7_EXP_PT_5_4_INV
    );
  EXP7_EXP_PT_5_5_INV_1469 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP7_EXP_PT_5_5_INV
    );
  EXP6_EXP_PT_0_0_INV_1470 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP6_EXP_PT_0_0_INV
    );
  EXP6_EXP_PT_0_2_INV_1471 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP6_EXP_PT_0_2_INV
    );
  EXP6_EXP_PT_0_3_INV_1472 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP6_EXP_PT_0_3_INV
    );
  EXP6_EXP_PT_0_4_INV_1473 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP6_EXP_PT_0_4_INV
    );
  EXP6_EXP_PT_0_5_INV_1474 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP6_EXP_PT_0_5_INV
    );
  EXP6_EXP_PT_0_6_INV_1475 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP6_EXP_PT_0_6_INV
    );
  EXP6_EXP_PT_1_0_INV_1476 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP6_EXP_PT_1_0_INV
    );
  EXP6_EXP_PT_1_1_INV_1477 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP6_EXP_PT_1_1_INV
    );
  EXP6_EXP_PT_1_2_INV_1478 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP6_EXP_PT_1_2_INV
    );
  EXP6_EXP_PT_1_3_INV_1479 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP6_EXP_PT_1_3_INV
    );
  EXP6_EXP_PT_1_4_INV_1480 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP6_EXP_PT_1_4_INV
    );
  EXP6_EXP_PT_1_5_INV_1481 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP6_EXP_PT_1_5_INV
    );
  EXP6_EXP_PT_2_1_INV_1482 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => EXP6_EXP_PT_2_1_INV
    );
  EXP6_EXP_PT_2_7_INV_1483 : X_INV 
    port map (
      I => LIGHT_VALUE(3),
      O => EXP6_EXP_PT_2_7_INV
    );
  EXP6_EXP_PT_2_8_INV_1484 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP6_EXP_PT_2_8_INV
    );
  EXP6_EXP_PT_3_1_INV_1485 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => EXP6_EXP_PT_3_1_INV
    );
  EXP6_EXP_PT_3_7_INV_1486 : X_INV 
    port map (
      I => LIGHT_VALUE(1),
      O => EXP6_EXP_PT_3_7_INV
    );
  EXP6_EXP_PT_3_8_INV_1487 : X_INV 
    port map (
      I => LIGHT_VALUE(2),
      O => EXP6_EXP_PT_3_8_INV
    );
  EXP6_EXP_PT_3_9_INV_1488 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP6_EXP_PT_3_9_INV
    );
  LIGHT_VALUE_3_SETF_PT_0_0_INV_1489 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => LIGHT_VALUE_3_SETF_PT_0_0_INV
    );
  LIGHT_VALUE_3_SETF_PT_0_1_INV_1490 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_3_SETF_PT_0_1_INV
    );
  LIGHT_VALUE_3_D2_PT_1_1_INV_1491 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_3_D2_PT_1_1_INV
    );
  LIGHT_VALUE_3_D2_PT_1_2_INV_1492 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_3_D2_PT_1_2_INV
    );
  LIGHT_VALUE_3_D2_PT_1_3_INV_1493 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => LIGHT_VALUE_3_D2_PT_1_3_INV
    );
  LIGHT_VALUE_3_D2_PT_1_4_INV_1494 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => LIGHT_VALUE_3_D2_PT_1_4_INV
    );
  LIGHT_VALUE_3_D2_PT_1_5_INV_1495 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => LIGHT_VALUE_3_D2_PT_1_5_INV
    );
  LIGHT_VALUE_3_D2_PT_1_6_INV_1496 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => LIGHT_VALUE_3_D2_PT_1_6_INV
    );
  LIGHT_VALUE_3_D2_PT_1_7_INV_1497 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => LIGHT_VALUE_3_D2_PT_1_7_INV
    );
  LIGHT_VALUE_3_D2_PT_1_8_INV_1498 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => LIGHT_VALUE_3_D2_PT_1_8_INV
    );
  LIGHT_VALUE_3_D2_PT_1_9_INV_1499 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => LIGHT_VALUE_3_D2_PT_1_9_INV
    );
  LIGHT_VALUE_3_D2_PT_1_10_INV_1500 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => LIGHT_VALUE_3_D2_PT_1_10_INV
    );
  LIGHT_VALUE_3_D2_PT_1_11_INV_1501 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => LIGHT_VALUE_3_D2_PT_1_11_INV
    );
  LIGHT_VALUE_3_D2_PT_1_12_INV_1502 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => LIGHT_VALUE_3_D2_PT_1_12_INV
    );
  LIGHT_VALUE_3_D2_PT_2_0_INV_1503 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => LIGHT_VALUE_3_D2_PT_2_0_INV
    );
  LIGHT_VALUE_3_D2_PT_2_2_INV_1504 : X_INV 
    port map (
      I => LIGHT_VALUE_5_FBK,
      O => LIGHT_VALUE_3_D2_PT_2_2_INV
    );
  LIGHT_VALUE_3_EXP_PT_0_1_INV_1505 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_3_EXP_PT_0_1_INV
    );
  LIGHT_VALUE_3_EXP_PT_0_3_INV_1506 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_3_EXP_PT_0_3_INV
    );
  LIGHT_VALUE_3_EXP_PT_0_4_INV_1507 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => LIGHT_VALUE_3_EXP_PT_0_4_INV
    );
  LIGHT_VALUE_3_EXP_PT_0_5_INV_1508 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => LIGHT_VALUE_3_EXP_PT_0_5_INV
    );
  LIGHT_VALUE_3_EXP_PT_0_6_INV_1509 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => LIGHT_VALUE_3_EXP_PT_0_6_INV
    );
  LIGHT_VALUE_3_EXP_PT_0_7_INV_1510 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => LIGHT_VALUE_3_EXP_PT_0_7_INV
    );
  LIGHT_VALUE_3_EXP_PT_0_8_INV_1511 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => LIGHT_VALUE_3_EXP_PT_0_8_INV
    );
  LIGHT_VALUE_3_EXP_PT_0_9_INV_1512 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => LIGHT_VALUE_3_EXP_PT_0_9_INV
    );
  LIGHT_VALUE_3_EXP_PT_0_10_INV_1513 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => LIGHT_VALUE_3_EXP_PT_0_10_INV
    );
  LIGHT_VALUE_3_EXP_PT_0_11_INV_1514 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => LIGHT_VALUE_3_EXP_PT_0_11_INV
    );
  LIGHT_VALUE_3_EXP_PT_0_12_INV_1515 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => LIGHT_VALUE_3_EXP_PT_0_12_INV
    );
  LIGHT_VALUE_3_EXP_PT_1_0_INV_1516 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => LIGHT_VALUE_3_EXP_PT_1_0_INV
    );
  LIGHT_VALUE_3_EXP_PT_1_12_INV_1517 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => LIGHT_VALUE_3_EXP_PT_1_12_INV
    );
  LIGHT_VALUE_3_EXP_PT_1_13_INV_1518 : X_INV 
    port map (
      I => LIGHT_VALUE(4),
      O => LIGHT_VALUE_3_EXP_PT_1_13_INV
    );
  FC1_CNT_6_RSTF_PT_0_0_INV_1519 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_6_RSTF_PT_0_0_INV
    );
  FC1_CNT_6_RSTF_PT_0_1_INV_1520 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_6_RSTF_PT_0_1_INV
    );
  FC1_CNT_6_D2_PT_2_7_INV_1521 : X_INV 
    port map (
      I => LIGHT_VALUE(5),
      O => FC1_CNT_6_D2_PT_2_7_INV
    );
  FC1_CNT_6_D2_PT_2_8_INV_1522 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => FC1_CNT_6_D2_PT_2_8_INV
    );
  FC1_CNT_6_D2_PT_3_0_INV_1523 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_6_D2_PT_3_0_INV
    );
  FC1_CNT_6_D2_PT_3_1_INV_1524 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => FC1_CNT_6_D2_PT_3_1_INV
    );
  FC1_CNT_6_D2_PT_3_2_INV_1525 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => FC1_CNT_6_D2_PT_3_2_INV
    );
  FC1_CNT_6_D2_PT_3_3_INV_1526 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => FC1_CNT_6_D2_PT_3_3_INV
    );
  FC1_CNT_6_D2_PT_3_4_INV_1527 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => FC1_CNT_6_D2_PT_3_4_INV
    );
  FC1_CNT_6_D2_PT_3_5_INV_1528 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => FC1_CNT_6_D2_PT_3_5_INV
    );
  FC1_CNT_6_D2_PT_3_7_INV_1529 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => FC1_CNT_6_D2_PT_3_7_INV
    );
  FC1_CNT_6_D2_PT_4_0_INV_1530 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_6_D2_PT_4_0_INV
    );
  FC1_CNT_6_D2_PT_4_1_INV_1531 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => FC1_CNT_6_D2_PT_4_1_INV
    );
  FC1_CNT_6_D2_PT_4_2_INV_1532 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => FC1_CNT_6_D2_PT_4_2_INV
    );
  FC1_CNT_6_D2_PT_4_3_INV_1533 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => FC1_CNT_6_D2_PT_4_3_INV
    );
  FC1_CNT_6_D2_PT_4_4_INV_1534 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => FC1_CNT_6_D2_PT_4_4_INV
    );
  FC1_CNT_6_D2_PT_4_5_INV_1535 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => FC1_CNT_6_D2_PT_4_5_INV
    );
  FC1_CNT_6_D2_PT_4_6_INV_1536 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => FC1_CNT_6_D2_PT_4_6_INV
    );
  FC1_CNT_6_D2_PT_5_0_INV_1537 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => FC1_CNT_6_D2_PT_5_0_INV
    );
  FC1_CNT_6_D2_PT_5_1_INV_1538 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => FC1_CNT_6_D2_PT_5_1_INV
    );
  FC1_CNT_6_D2_PT_5_2_INV_1539 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => FC1_CNT_6_D2_PT_5_2_INV
    );
  FC1_CNT_6_D2_PT_5_3_INV_1540 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => FC1_CNT_6_D2_PT_5_3_INV
    );
  FC1_CNT_6_D2_PT_5_4_INV_1541 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => FC1_CNT_6_D2_PT_5_4_INV
    );
  FC1_CNT_6_D2_PT_5_5_INV_1542 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => FC1_CNT_6_D2_PT_5_5_INV
    );
  FC1_CNT_6_D2_PT_5_6_INV_1543 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => FC1_CNT_6_D2_PT_5_6_INV
    );
  EXP5_EXP_PT_0_0_INV_1544 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP5_EXP_PT_0_0_INV
    );
  EXP5_EXP_PT_0_2_INV_1545 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP5_EXP_PT_0_2_INV
    );
  EXP5_EXP_PT_0_3_INV_1546 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP5_EXP_PT_0_3_INV
    );
  EXP5_EXP_PT_0_4_INV_1547 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP5_EXP_PT_0_4_INV
    );
  EXP5_EXP_PT_0_5_INV_1548 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP5_EXP_PT_0_5_INV
    );
  EXP5_EXP_PT_0_6_INV_1549 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => EXP5_EXP_PT_0_6_INV
    );
  EXP5_EXP_PT_0_7_INV_1550 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP5_EXP_PT_0_7_INV
    );
  EXP5_EXP_PT_1_0_INV_1551 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP5_EXP_PT_1_0_INV
    );
  EXP5_EXP_PT_1_1_INV_1552 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP5_EXP_PT_1_1_INV
    );
  EXP5_EXP_PT_1_2_INV_1553 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP5_EXP_PT_1_2_INV
    );
  EXP5_EXP_PT_1_3_INV_1554 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP5_EXP_PT_1_3_INV
    );
  EXP5_EXP_PT_1_4_INV_1555 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP5_EXP_PT_1_4_INV
    );
  EXP5_EXP_PT_1_5_INV_1556 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => EXP5_EXP_PT_1_5_INV
    );
  EXP5_EXP_PT_1_6_INV_1557 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP5_EXP_PT_1_6_INV
    );
  EXP5_EXP_PT_2_0_INV_1558 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_1_FBK,
      O => EXP5_EXP_PT_2_0_INV
    );
  EXP5_EXP_PT_2_1_INV_1559 : X_INV 
    port map (
      I => FC1_CNT_3_FBK,
      O => EXP5_EXP_PT_2_1_INV
    );
  EXP5_EXP_PT_2_2_INV_1560 : X_INV 
    port map (
      I => FC1_CNT(1),
      O => EXP5_EXP_PT_2_2_INV
    );
  EXP5_EXP_PT_2_3_INV_1561 : X_INV 
    port map (
      I => FC1_CNT(2),
      O => EXP5_EXP_PT_2_3_INV
    );
  EXP5_EXP_PT_2_4_INV_1562 : X_INV 
    port map (
      I => FC1_CNT_4_FBK,
      O => EXP5_EXP_PT_2_4_INV
    );
  EXP5_EXP_PT_2_5_INV_1563 : X_INV 
    port map (
      I => FC1_CNT_5_FBK,
      O => EXP5_EXP_PT_2_5_INV
    );
  EXP5_EXP_PT_2_6_INV_1564 : X_INV 
    port map (
      I => FC1_CNT(0),
      O => EXP5_EXP_PT_2_6_INV
    );
  EXP5_EXP_PT_3_1_INV_1565 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => EXP5_EXP_PT_3_1_INV
    );
  EXP5_EXP_PT_3_8_INV_1566 : X_INV 
    port map (
      I => LIGHT_VALUE(3),
      O => EXP5_EXP_PT_3_8_INV
    );
  EXP5_EXP_PT_3_9_INV_1567 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP5_EXP_PT_3_9_INV
    );
  EXP5_EXP_PT_4_1_INV_1568 : X_INV 
    port map (
      I => LIGHT_VALUE_4_FBK,
      O => EXP5_EXP_PT_4_1_INV
    );
  EXP5_EXP_PT_4_8_INV_1569 : X_INV 
    port map (
      I => LIGHT_VALUE(1),
      O => EXP5_EXP_PT_4_8_INV
    );
  EXP5_EXP_PT_4_9_INV_1570 : X_INV 
    port map (
      I => LIGHT_VALUE(2),
      O => EXP5_EXP_PT_4_9_INV
    );
  EXP5_EXP_PT_4_10_INV_1571 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE_0_FBK,
      O => EXP5_EXP_PT_4_10_INV
    );
  LIGHT_VALUE_0_RSTF_PT_0_0_INV_1572 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => LIGHT_VALUE_0_RSTF_PT_0_0_INV
    );
  LIGHT_VALUE_0_RSTF_PT_0_1_INV_1573 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_0_RSTF_PT_0_1_INV
    );
  LIGHT_VALUE_0_D2_PT_2_1_INV_1574 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_0_D2_PT_2_1_INV
    );
  LIGHT_VALUE_0_D2_PT_2_2_INV_1575 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_0_D2_PT_2_2_INV
    );
  LIGHT_VALUE_0_D2_PT_2_3_INV_1576 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => LIGHT_VALUE_0_D2_PT_2_3_INV
    );
  LIGHT_VALUE_0_D2_PT_2_4_INV_1577 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => LIGHT_VALUE_0_D2_PT_2_4_INV
    );
  LIGHT_VALUE_0_D2_PT_2_5_INV_1578 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => LIGHT_VALUE_0_D2_PT_2_5_INV
    );
  LIGHT_VALUE_0_D2_PT_2_6_INV_1579 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => LIGHT_VALUE_0_D2_PT_2_6_INV
    );
  LIGHT_VALUE_0_D2_PT_2_7_INV_1580 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => LIGHT_VALUE_0_D2_PT_2_7_INV
    );
  LIGHT_VALUE_0_D2_PT_2_8_INV_1581 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => LIGHT_VALUE_0_D2_PT_2_8_INV
    );
  LIGHT_VALUE_0_D2_PT_2_9_INV_1582 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => LIGHT_VALUE_0_D2_PT_2_9_INV
    );
  LIGHT_VALUE_0_D2_PT_3_1_INV_1583 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_0_D2_PT_3_1_INV
    );
  LIGHT_VALUE_0_D2_PT_3_2_INV_1584 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_0_D2_PT_3_2_INV
    );
  LIGHT_VALUE_0_D2_PT_3_3_INV_1585 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => LIGHT_VALUE_0_D2_PT_3_3_INV
    );
  LIGHT_VALUE_0_D2_PT_3_4_INV_1586 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => LIGHT_VALUE_0_D2_PT_3_4_INV
    );
  LIGHT_VALUE_0_D2_PT_3_5_INV_1587 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => LIGHT_VALUE_0_D2_PT_3_5_INV
    );
  LIGHT_VALUE_0_D2_PT_3_6_INV_1588 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => LIGHT_VALUE_0_D2_PT_3_6_INV
    );
  LIGHT_VALUE_0_D2_PT_3_7_INV_1589 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => LIGHT_VALUE_0_D2_PT_3_7_INV
    );
  LIGHT_VALUE_0_D2_PT_3_8_INV_1590 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => LIGHT_VALUE_0_D2_PT_3_8_INV
    );
  LIGHT_VALUE_0_D2_PT_3_9_INV_1591 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => LIGHT_VALUE_0_D2_PT_3_9_INV
    );
  LIGHT_VALUE_0_D2_PT_4_1_INV_1592 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_0_D2_PT_4_1_INV
    );
  LIGHT_VALUE_0_D2_PT_4_2_INV_1593 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_0_D2_PT_4_2_INV
    );
  LIGHT_VALUE_0_D2_PT_4_3_INV_1594 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => LIGHT_VALUE_0_D2_PT_4_3_INV
    );
  LIGHT_VALUE_0_D2_PT_4_4_INV_1595 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => LIGHT_VALUE_0_D2_PT_4_4_INV
    );
  LIGHT_VALUE_0_D2_PT_4_5_INV_1596 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => LIGHT_VALUE_0_D2_PT_4_5_INV
    );
  LIGHT_VALUE_0_D2_PT_4_6_INV_1597 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => LIGHT_VALUE_0_D2_PT_4_6_INV
    );
  LIGHT_VALUE_0_D2_PT_4_7_INV_1598 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => LIGHT_VALUE_0_D2_PT_4_7_INV
    );
  LIGHT_VALUE_0_D2_PT_4_8_INV_1599 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => LIGHT_VALUE_0_D2_PT_4_8_INV
    );
  LIGHT_VALUE_0_D2_PT_4_9_INV_1600 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => LIGHT_VALUE_0_D2_PT_4_9_INV
    );
  LIGHT_VALUE_0_D2_PT_5_0_INV_1601 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => LIGHT_VALUE_0_D2_PT_5_0_INV
    );
  LIGHT_VALUE_0_D2_PT_5_2_INV_1602 : X_INV 
    port map (
      I => LIGHT_VALUE_5_FBK,
      O => LIGHT_VALUE_0_D2_PT_5_2_INV
    );
  TD1_CNT_5_SETF_PT_0_0_INV_1603 : X_INV 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM,
      O => TD1_CNT_5_SETF_PT_0_0_INV
    );
  TD1_CNT_5_SETF_PT_0_1_INV_1604 : X_INV 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM,
      O => TD1_CNT_5_SETF_PT_0_1_INV
    );
  TD1_CNT_5_D2_PT_0_0_INV_1605 : X_INV 
    port map (
      I => TD1_CNT_0_FBK,
      O => TD1_CNT_5_D2_PT_0_0_INV
    );
  TD1_CNT_5_D2_PT_0_1_INV_1606 : X_INV 
    port map (
      I => TD1_CNT_1_Q_3,
      O => TD1_CNT_5_D2_PT_0_1_INV
    );
  TD1_CNT_5_D2_PT_0_2_INV_1607 : X_INV 
    port map (
      I => TD1_CNT_2_FBK,
      O => TD1_CNT_5_D2_PT_0_2_INV
    );
  TD1_CNT_5_D2_PT_0_3_INV_1608 : X_INV 
    port map (
      I => TD1_CNT_3_FBK,
      O => TD1_CNT_5_D2_PT_0_3_INV
    );
  TD1_CNT_5_D2_PT_0_4_INV_1609 : X_INV 
    port map (
      I => TD1_CNT_4_FBK,
      O => TD1_CNT_5_D2_PT_0_4_INV
    );
  TD1_CNT_5_EXP_PT_0_1_INV_1610 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => TD1_CNT_5_EXP_PT_0_1_INV
    );
  TD1_CNT_5_EXP_PT_0_3_INV_1611 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => TD1_CNT_5_EXP_PT_0_3_INV
    );
  TD1_CNT_5_EXP_PT_0_4_INV_1612 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => TD1_CNT_5_EXP_PT_0_4_INV
    );
  TD1_CNT_5_EXP_PT_0_5_INV_1613 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => TD1_CNT_5_EXP_PT_0_5_INV
    );
  TD1_CNT_5_EXP_PT_0_6_INV_1614 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => TD1_CNT_5_EXP_PT_0_6_INV
    );
  TD1_CNT_5_EXP_PT_0_7_INV_1615 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => TD1_CNT_5_EXP_PT_0_7_INV
    );
  TD1_CNT_5_EXP_PT_0_8_INV_1616 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => TD1_CNT_5_EXP_PT_0_8_INV
    );
  TD1_CNT_5_EXP_PT_0_9_INV_1617 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => TD1_CNT_5_EXP_PT_0_9_INV
    );
  TD1_CNT_5_EXP_PT_0_10_INV_1618 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => TD1_CNT_5_EXP_PT_0_10_INV
    );
  TD1_CNT_5_EXP_PT_1_0_INV_1619 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => TD1_CNT_5_EXP_PT_1_0_INV
    );
  TD1_CNT_5_EXP_PT_1_10_INV_1620 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => TD1_CNT_5_EXP_PT_1_10_INV
    );
  TD1_CNT_5_EXP_PT_1_11_INV_1621 : X_INV 
    port map (
      I => LIGHT_VALUE(4),
      O => TD1_CNT_5_EXP_PT_1_11_INV
    );
  TD1_CNT_5_EXP_PT_2_0_INV_1622 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => TD1_CNT_5_EXP_PT_2_0_INV
    );
  TD1_CNT_5_EXP_PT_2_10_INV_1623 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => TD1_CNT_5_EXP_PT_2_10_INV
    );
  TD1_CNT_5_EXP_PT_2_11_INV_1624 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => TD1_CNT_5_EXP_PT_2_11_INV
    );
  TD1_CNT_5_EXP_PT_2_12_INV_1625 : X_INV 
    port map (
      I => LIGHT_VALUE(4),
      O => TD1_CNT_5_EXP_PT_2_12_INV
    );
  TD1_CNT_1_SETF_PT_0_0_INV_1626 : X_INV 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_FBK,
      O => TD1_CNT_1_SETF_PT_0_0_INV
    );
  TD1_CNT_1_SETF_PT_0_1_INV_1627 : X_INV 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_FBK,
      O => TD1_CNT_1_SETF_PT_0_1_INV
    );
  TD1_CNT_1_XOR_0_INV_1628 : X_INV 
    port map (
      I => TD1_CNT_1_D1,
      O => TD1_CNT_1_XOR_0_INV
    );
  TD1_CNT_2_RSTF_PT_0_0_INV_1629 : X_INV 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM,
      O => TD1_CNT_2_RSTF_PT_0_0_INV
    );
  TD1_CNT_2_RSTF_PT_0_1_INV_1630 : X_INV 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM,
      O => TD1_CNT_2_RSTF_PT_0_1_INV
    );
  TD1_CNT_2_D2_PT_0_0_INV_1631 : X_INV 
    port map (
      I => TD1_CNT_0_FBK,
      O => TD1_CNT_2_D2_PT_0_0_INV
    );
  TD1_CNT_2_D2_PT_0_1_INV_1632 : X_INV 
    port map (
      I => TD1_CNT_1_Q_3,
      O => TD1_CNT_2_D2_PT_0_1_INV
    );
  TD1_CNT_3_EXP_PT_0_0_INV_1633 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => TD1_CNT_3_EXP_PT_0_0_INV
    );
  TD1_CNT_3_EXP_PT_0_1_INV_1634 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => TD1_CNT_3_EXP_PT_0_1_INV
    );
  TD1_CNT_3_EXP_PT_0_2_INV_1635 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => TD1_CNT_3_EXP_PT_0_2_INV
    );
  TD1_CNT_3_EXP_PT_0_3_INV_1636 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => TD1_CNT_3_EXP_PT_0_3_INV
    );
  TD1_CNT_3_EXP_PT_1_0_INV_1637 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => TD1_CNT_3_EXP_PT_1_0_INV
    );
  TD1_CNT_3_EXP_PT_1_1_INV_1638 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => TD1_CNT_3_EXP_PT_1_1_INV
    );
  TD1_CNT_3_EXP_PT_1_2_INV_1639 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => TD1_CNT_3_EXP_PT_1_2_INV
    );
  TD1_CNT_3_SETF_PT_0_0_INV_1640 : X_INV 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM,
      O => TD1_CNT_3_SETF_PT_0_0_INV
    );
  TD1_CNT_3_SETF_PT_0_1_INV_1641 : X_INV 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM,
      O => TD1_CNT_3_SETF_PT_0_1_INV
    );
  TD1_CNT_3_D2_PT_0_0_INV_1642 : X_INV 
    port map (
      I => TD1_CNT_0_FBK,
      O => TD1_CNT_3_D2_PT_0_0_INV
    );
  TD1_CNT_3_D2_PT_0_1_INV_1643 : X_INV 
    port map (
      I => TD1_CNT_1_Q_3,
      O => TD1_CNT_3_D2_PT_0_1_INV
    );
  TD1_CNT_3_D2_PT_0_2_INV_1644 : X_INV 
    port map (
      I => TD1_CNT_2_FBK,
      O => TD1_CNT_3_D2_PT_0_2_INV
    );
  LIGHT_VALUE_2_RSTF_PT_0_0_INV_1645 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => LIGHT_VALUE_2_RSTF_PT_0_0_INV
    );
  LIGHT_VALUE_2_RSTF_PT_0_1_INV_1646 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_2_RSTF_PT_0_1_INV
    );
  LIGHT_VALUE_2_D2_PT_1_1_INV_1647 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_2_D2_PT_1_1_INV
    );
  LIGHT_VALUE_2_D2_PT_1_2_INV_1648 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_2_D2_PT_1_2_INV
    );
  LIGHT_VALUE_2_D2_PT_1_3_INV_1649 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => LIGHT_VALUE_2_D2_PT_1_3_INV
    );
  LIGHT_VALUE_2_D2_PT_1_4_INV_1650 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => LIGHT_VALUE_2_D2_PT_1_4_INV
    );
  LIGHT_VALUE_2_D2_PT_1_5_INV_1651 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => LIGHT_VALUE_2_D2_PT_1_5_INV
    );
  LIGHT_VALUE_2_D2_PT_1_6_INV_1652 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => LIGHT_VALUE_2_D2_PT_1_6_INV
    );
  LIGHT_VALUE_2_D2_PT_1_7_INV_1653 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => LIGHT_VALUE_2_D2_PT_1_7_INV
    );
  LIGHT_VALUE_2_D2_PT_1_8_INV_1654 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => LIGHT_VALUE_2_D2_PT_1_8_INV
    );
  LIGHT_VALUE_2_D2_PT_1_9_INV_1655 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => LIGHT_VALUE_2_D2_PT_1_9_INV
    );
  LIGHT_VALUE_2_D2_PT_1_10_INV_1656 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => LIGHT_VALUE_2_D2_PT_1_10_INV
    );
  LIGHT_VALUE_2_D2_PT_1_12_INV_1657 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => LIGHT_VALUE_2_D2_PT_1_12_INV
    );
  LIGHT_VALUE_2_D2_PT_2_1_INV_1658 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_2_D2_PT_2_1_INV
    );
  LIGHT_VALUE_2_D2_PT_2_2_INV_1659 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_2_D2_PT_2_2_INV
    );
  LIGHT_VALUE_2_D2_PT_2_3_INV_1660 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => LIGHT_VALUE_2_D2_PT_2_3_INV
    );
  LIGHT_VALUE_2_D2_PT_2_4_INV_1661 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => LIGHT_VALUE_2_D2_PT_2_4_INV
    );
  LIGHT_VALUE_2_D2_PT_2_5_INV_1662 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => LIGHT_VALUE_2_D2_PT_2_5_INV
    );
  LIGHT_VALUE_2_D2_PT_2_6_INV_1663 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => LIGHT_VALUE_2_D2_PT_2_6_INV
    );
  LIGHT_VALUE_2_D2_PT_2_7_INV_1664 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => LIGHT_VALUE_2_D2_PT_2_7_INV
    );
  LIGHT_VALUE_2_D2_PT_2_8_INV_1665 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => LIGHT_VALUE_2_D2_PT_2_8_INV
    );
  LIGHT_VALUE_2_D2_PT_2_9_INV_1666 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => LIGHT_VALUE_2_D2_PT_2_9_INV
    );
  LIGHT_VALUE_2_D2_PT_2_10_INV_1667 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => LIGHT_VALUE_2_D2_PT_2_10_INV
    );
  LIGHT_VALUE_2_D2_PT_2_11_INV_1668 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => LIGHT_VALUE_2_D2_PT_2_11_INV
    );
  LIGHT_VALUE_2_D2_PT_3_1_INV_1669 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(1),
      O => LIGHT_VALUE_2_D2_PT_3_1_INV
    );
  LIGHT_VALUE_2_D2_PT_3_2_INV_1670 : X_INV 
    port map (
      I => FC1_CNT_1_FBK,
      O => LIGHT_VALUE_2_D2_PT_3_2_INV
    );
  LIGHT_VALUE_2_D2_PT_3_3_INV_1671 : X_INV 
    port map (
      I => FC1_CNT_2_FBK,
      O => LIGHT_VALUE_2_D2_PT_3_3_INV
    );
  LIGHT_VALUE_2_D2_PT_3_4_INV_1672 : X_INV 
    port map (
      I => FC1_CNT_0_FBK,
      O => LIGHT_VALUE_2_D2_PT_3_4_INV
    );
  LIGHT_VALUE_2_D2_PT_3_5_INV_1673 : X_INV 
    port map (
      I => FC1_CNT(3),
      O => LIGHT_VALUE_2_D2_PT_3_5_INV
    );
  LIGHT_VALUE_2_D2_PT_3_6_INV_1674 : X_INV 
    port map (
      I => FC1_CNT(4),
      O => LIGHT_VALUE_2_D2_PT_3_6_INV
    );
  LIGHT_VALUE_2_D2_PT_3_7_INV_1675 : X_INV 
    port map (
      I => FC1_CNT(5),
      O => LIGHT_VALUE_2_D2_PT_3_7_INV
    );
  LIGHT_VALUE_2_D2_PT_3_8_INV_1676 : X_INV 
    port map (
      I => FC1_CNT(6),
      O => LIGHT_VALUE_2_D2_PT_3_8_INV
    );
  LIGHT_VALUE_2_D2_PT_3_9_INV_1677 : X_INV 
    port map (
      I => FC1_CNT(7),
      O => LIGHT_VALUE_2_D2_PT_3_9_INV
    );
  LIGHT_VALUE_2_D2_PT_3_10_INV_1678 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => LIGHT_VALUE_2_D2_PT_3_10_INV
    );
  LIGHT_VALUE_2_D2_PT_3_11_INV_1679 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => LIGHT_VALUE_2_D2_PT_3_11_INV
    );
  LIGHT_VALUE_2_D2_PT_4_0_INV_1680 : X_INV 
    port map (
      I => DFSM1_CURRENT_STATE_H_CURRENT_STATE(0),
      O => LIGHT_VALUE_2_D2_PT_4_0_INV
    );
  LIGHT_VALUE_2_D2_PT_4_2_INV_1681 : X_INV 
    port map (
      I => LIGHT_VALUE_5_FBK,
      O => LIGHT_VALUE_2_D2_PT_4_2_INV
    );
  TD1_CNT_4_RSTF_PT_0_0_INV_1682 : X_INV 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM,
      O => TD1_CNT_4_RSTF_PT_0_0_INV
    );
  TD1_CNT_4_RSTF_PT_0_1_INV_1683 : X_INV 
    port map (
      I => TD1_CNT_5_TD1_CNT_5_SETF_INT_UIM,
      O => TD1_CNT_4_RSTF_PT_0_1_INV
    );
  TD1_CNT_4_D2_PT_0_0_INV_1684 : X_INV 
    port map (
      I => TD1_CNT_0_FBK,
      O => TD1_CNT_4_D2_PT_0_0_INV
    );
  TD1_CNT_4_D2_PT_0_1_INV_1685 : X_INV 
    port map (
      I => TD1_CNT_1_Q_3,
      O => TD1_CNT_4_D2_PT_0_1_INV
    );
  TD1_CNT_4_D2_PT_0_2_INV_1686 : X_INV 
    port map (
      I => TD1_CNT_2_FBK,
      O => TD1_CNT_4_D2_PT_0_2_INV
    );
  TD1_CNT_4_D2_PT_0_3_INV_1687 : X_INV 
    port map (
      I => TD1_CNT_3_FBK,
      O => TD1_CNT_4_D2_PT_0_3_INV
    );
  TD1_CNT_4_EXP_PT_0_0_INV_1688 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => TD1_CNT_4_EXP_PT_0_0_INV
    );
  TD1_CNT_4_EXP_PT_0_1_INV_1689 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => TD1_CNT_4_EXP_PT_0_1_INV
    );
  TD1_CNT_4_EXP_PT_0_2_INV_1690 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => TD1_CNT_4_EXP_PT_0_2_INV
    );
  TD1_CNT_4_EXP_PT_1_0_INV_1691 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => TD1_CNT_4_EXP_PT_1_0_INV
    );
  TD1_CNT_4_EXP_PT_1_1_INV_1692 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => TD1_CNT_4_EXP_PT_1_1_INV
    );
  TD1_CNT_4_EXP_PT_2_0_INV_1693 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => TD1_CNT_4_EXP_PT_2_0_INV
    );
  CM_FADE_UP_D2_PT_2_0_INV_1694 : X_INV 
    port map (
      I => RXD_READY_FBK,
      O => CM_FADE_UP_D2_PT_2_0_INV
    );
  CM_FADE_UP_D2_PT_2_1_INV_1695 : X_INV 
    port map (
      I => RXD_READY_FBK,
      O => CM_FADE_UP_D2_PT_2_1_INV
    );
  CM_FADE_UP_D2_PT_5_1_INV_1696 : X_INV 
    port map (
      I => RXD_4_FBK,
      O => CM_FADE_UP_D2_PT_5_1_INV
    );
  CM_FADE_UP_D2_PT_6_0_INV_1697 : X_INV 
    port map (
      I => RC_ADDRESS_C(0),
      O => CM_FADE_UP_D2_PT_6_0_INV
    );
  CM_FADE_UP_XOR_0_INV_1698 : X_INV 
    port map (
      I => CM_FADE_UP_D1,
      O => CM_FADE_UP_XOR_0_INV
    );
  EXP15_EXP_PT_1_1_INV_1699 : X_INV 
    port map (
      I => CM_FADE_UP_FBK,
      O => EXP15_EXP_PT_1_1_INV
    );
  EXP15_EXP_PT_3_0_INV_1700 : X_INV 
    port map (
      I => RXD_1_FBK,
      O => EXP15_EXP_PT_3_0_INV
    );
  EXP15_EXP_PT_3_1_INV_1701 : X_INV 
    port map (
      I => CM_FADE_UP_FBK,
      O => EXP15_EXP_PT_3_1_INV
    );
  EXP15_EXP_PT_4_1_INV_1702 : X_INV 
    port map (
      I => CM_FADE_UP_FBK,
      O => EXP15_EXP_PT_4_1_INV
    );
  EXP15_EXP_PT_5_0_INV_1703 : X_INV 
    port map (
      I => RC_ADDRESS_C(3),
      O => EXP15_EXP_PT_5_0_INV
    );
  EXP16_EXP_PT_1_0_INV_1704 : X_INV 
    port map (
      I => RXD_3_FBK,
      O => EXP16_EXP_PT_1_0_INV
    );
  EXP16_EXP_PT_1_1_INV_1705 : X_INV 
    port map (
      I => RXD_0_FBK,
      O => EXP16_EXP_PT_1_1_INV
    );
  Q_OPTX_FX_DC_68_D2_PT_2_0_INV_1706 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => Q_OPTX_FX_DC_68_D2_PT_2_0_INV
    );
  Q_OPTX_FX_DC_68_D2_PT_3_0_INV_1707 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => Q_OPTX_FX_DC_68_D2_PT_3_0_INV
    );
  Q_OPTX_FX_DC_68_D2_PT_3_1_INV_1708 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => Q_OPTX_FX_DC_68_D2_PT_3_1_INV
    );
  Q_OPTX_FX_DC_68_D2_PT_4_0_INV_1709 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => Q_OPTX_FX_DC_68_D2_PT_4_0_INV
    );
  Q_OPTX_FX_DC_68_D2_PT_5_0_INV_1710 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => Q_OPTX_FX_DC_68_D2_PT_5_0_INV
    );
  Q_OPTX_FX_DC_68_D2_PT_5_1_INV_1711 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => Q_OPTX_FX_DC_68_D2_PT_5_1_INV
    );
  Q_OPTX_FX_DC_68_D2_PT_6_0_INV_1712 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => Q_OPTX_FX_DC_68_D2_PT_6_0_INV
    );
  EXP11_EXP_PT_1_0_INV_1713 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => EXP11_EXP_PT_1_0_INV
    );
  EXP11_EXP_PT_1_1_INV_1714 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => EXP11_EXP_PT_1_1_INV
    );
  EXP11_EXP_PT_1_2_INV_1715 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => EXP11_EXP_PT_1_2_INV
    );
  EXP11_EXP_PT_2_0_INV_1716 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => EXP11_EXP_PT_2_0_INV
    );
  EXP11_EXP_PT_2_1_INV_1717 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => EXP11_EXP_PT_2_1_INV
    );
  EXP11_EXP_PT_2_2_INV_1718 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => EXP11_EXP_PT_2_2_INV
    );
  EXP11_EXP_PT_3_0_INV_1719 : X_INV 
    port map (
      I => LIGHT_VALUE_1_FBK,
      O => EXP11_EXP_PT_3_0_INV
    );
  EXP11_EXP_PT_3_1_INV_1720 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => EXP11_EXP_PT_3_1_INV
    );
  EXP11_EXP_PT_4_0_INV_1721 : X_INV 
    port map (
      I => LIGHT_VALUE_2_FBK,
      O => EXP11_EXP_PT_4_0_INV
    );
  EXP11_EXP_PT_4_1_INV_1722 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => EXP11_EXP_PT_4_1_INV
    );
  EXP11_EXP_PT_5_0_INV_1723 : X_INV 
    port map (
      I => LIGHT_VALUE_0_FBK,
      O => EXP11_EXP_PT_5_0_INV
    );
  EXP11_EXP_PT_5_1_INV_1724 : X_INV 
    port map (
      I => LIGHT_VALUE_3_FBK,
      O => EXP11_EXP_PT_5_1_INV
    );
  ROC_NGD2VHDL : ROC port map (O => PRLD);
end STRUCTURE;

